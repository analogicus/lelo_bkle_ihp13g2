magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747899951
<< checkpaint >>
rect 0 0 1 1
<< metal1 >>
rect -100 3930 5786 3980
<< metal1 >>
rect -100 -100 5786 -50
<< metal2 >>
rect -100 -50 -50 3930
<< metal2 >>
rect 5736 -50 5786 3930
<< metal1 >>
rect -107 3923 -43 3987
<< metal2 >>
rect -107 3923 -43 3987
<< via1 >>
rect -100 3930 -50 3980
<< metal1 >>
rect -107 -107 -43 -43
<< metal2 >>
rect -107 -107 -43 -43
<< via1 >>
rect -100 -100 -50 -50
<< metal1 >>
rect 5729 3923 5793 3987
<< metal2 >>
rect 5729 3923 5793 3987
<< via1 >>
rect 5736 3930 5786 3980
<< metal1 >>
rect 5729 -107 5793 -43
<< metal2 >>
rect 5729 -107 5793 -43
<< via1 >>
rect 5736 -100 5786 -50
<< metal1 >>
rect -200 4030 5886 4080
<< metal1 >>
rect -200 -200 5886 -150
<< metal2 >>
rect -200 -150 -150 4030
<< metal2 >>
rect 5836 -150 5886 4030
<< metal1 >>
rect -207 4023 -143 4087
<< metal2 >>
rect -207 4023 -143 4087
<< via1 >>
rect -200 4030 -150 4080
<< metal1 >>
rect -207 -207 -143 -143
<< metal2 >>
rect -207 -207 -143 -143
<< via1 >>
rect -200 -200 -150 -150
<< metal1 >>
rect 5829 4023 5893 4087
<< metal2 >>
rect 5829 4023 5893 4087
<< via1 >>
rect 5836 4030 5886 4080
<< metal1 >>
rect 5829 -207 5893 -143
<< metal2 >>
rect 5829 -207 5893 -143
<< via1 >>
rect 5836 -200 5886 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 5736 3930
<< labels >>
flabel metal1 s -200 4030 5886 4080 0 FreeSans 400 0 0 0 VDD_1V8
port 53 nsew signal bidirectional
flabel metal1 s -100 3930 5786 3980 0 FreeSans 400 0 0 0 VSS
port 54 nsew signal bidirectional
<< properties >>
<< end >>