magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747899951
<< checkpaint >>
rect 0 0 1 1
use LELOATR_PCH_4C5F0  diff1_MP3<3> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 964
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP3<2> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 964
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP3<1> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 1764
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  diff1_MP3<1>_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 2164
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP3<0> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 1764
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  diff1_MP3<0>_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 2164
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<3> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 2264
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  diff1_MP4<3>_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 2664
box 0 0 756 240
use LELOATR_PCH_4CTAPBOT  diff1_MP4<3>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 2024
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<2> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 2264
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  diff1_MP4<2>_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 2664
box 0 0 756 240
use LELOATR_PCH_4CTAPBOT  diff1_MP4<2>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 2024
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<1> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 564
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  diff1_MP4<1>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 324
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<0> ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 564
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  diff1_MP4<0>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 324
box 0 0 756 240
use LELOATR_PCH_4C5F0  mirror1_MP2 ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 1364
box 0 0 756 400
use LELOATR_PCH_4C5F0  mirror1_MP1 ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 1364
box 0 0 756 400
use LELOATR_NCH_4C5F0  mirror2_MN1 ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 3280
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN1_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 3680
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror2_MN1_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 1082 0 1 3040
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN2 ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 3280
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN2_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 3680
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror2_MN2_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747899951
transform 1 0 326 0 1 3040
box 0 0 756 240
use LELOTR_RPPO16  bias1_RH1 ../LELO_TR_IHP13G2
timestamp 1747899951
transform 1 0 2038 0 1 200
box 0 0 3448 880
use LELOTR_RPPO16  bias1_RH2 ../LELO_TR_IHP13G2
timestamp 1747899951
transform 1 0 2038 0 1 2060
box 0 0 3448 880
use LELOTR_RPPO16  bias1_RH3 ../LELO_TR_IHP13G2
timestamp 1747899951
transform 1 0 2038 0 1 1130
box 0 0 3448 880
<< metal3 >>
rect 454 1947 1221 1977
<< metal3 >>
rect 1063 1947 1221 1977
<< metal4 >>
rect 1063 1147 1093 1977
<< metal3 >>
rect 1063 1147 1221 1177
<< metal3 >>
rect 454 1147 1221 1177
<< metal3 >>
rect 1056 1940 1100 1984
<< metal4 >>
rect 1056 1940 1100 1984
<< via3 >>
rect 1063 1947 1093 1977
<< metal3 >>
rect 1056 1140 1100 1184
<< metal4 >>
rect 1056 1140 1100 1184
<< via3 >>
rect 1063 1147 1093 1177
<< metal3 >>
rect 439 749 1206 779
<< metal3 >>
rect 311 749 469 779
<< metal4 >>
rect 311 749 341 2475
<< metal3 >>
rect 311 2445 469 2475
<< metal3 >>
rect 439 2445 1206 2475
<< metal3 >>
rect 304 742 348 786
<< metal4 >>
rect 304 742 348 786
<< via3 >>
rect 311 749 341 779
<< metal3 >>
rect 304 2438 348 2482
<< metal4 >>
rect 304 2438 348 2482
<< via3 >>
rect 311 2445 341 2475
<< metal4 >>
rect 808 2285 838 3324
<< metal3 >>
rect 808 2285 1606 2315
<< metal3 >>
rect 1576 2285 1750 2315
<< metal4 >>
rect 1720 589 1750 2315
<< metal3 >>
rect 1576 589 1750 619
<< metal3 >>
rect 823 589 1606 619
<< metal3 >>
rect 801 2278 845 2322
<< metal4 >>
rect 801 2278 845 2322
<< via3 >>
rect 808 2285 838 2315
<< metal3 >>
rect 1713 2278 1757 2322
<< metal4 >>
rect 1713 2278 1757 2322
<< via3 >>
rect 1720 2285 1750 2315
<< metal3 >>
rect 1713 582 1757 626
<< metal4 >>
rect 1713 582 1757 626
<< via3 >>
rect 1720 589 1750 619
<< metal3 >>
rect 440 3467 1207 3497
<< metal3 >>
rect 440 3467 982 3497
<< metal4 >>
rect 952 1787 982 3497
<< metal3 >>
rect 808 1787 982 1817
<< metal3 >>
rect 808 1787 1606 1817
<< metal3 >>
rect 1576 1787 1846 1817
<< metal4 >>
rect 1816 987 1846 1817
<< metal3 >>
rect 1576 987 1846 1017
<< metal3 >>
rect 823 987 1606 1017
<< metal3 >>
rect 945 3460 989 3504
<< metal4 >>
rect 945 3460 989 3504
<< via3 >>
rect 952 3467 982 3497
<< metal3 >>
rect 945 1780 989 1824
<< metal4 >>
rect 945 1780 989 1824
<< via3 >>
rect 952 1787 982 1817
<< metal3 >>
rect 1809 1780 1853 1824
<< metal4 >>
rect 1809 1780 1853 1824
<< via3 >>
rect 1816 1787 1846 1817
<< metal3 >>
rect 1809 980 1853 1024
<< metal4 >>
rect 1809 980 1853 1024
<< via3 >>
rect 1816 987 1846 1017
<< metal3 >>
rect 1317 1382 1588 1412
<< metal4 >>
rect 1317 870 1347 1412
<< metal4 >>
rect 1317 870 1347 1300
<< metal3 >>
rect 1317 1270 1939 1300
<< metal4 >>
rect 1909 1270 1939 2100
<< metal3 >>
rect 1317 2070 1939 2100
<< metal4 >>
rect 1317 2070 1347 2596
<< metal3 >>
rect 565 2566 1347 2596
<< metal4 >>
rect 565 2070 595 2596
<< metal3 >>
rect 213 2070 595 2100
<< metal4 >>
rect 213 1270 243 2100
<< metal3 >>
rect 213 1270 595 1300
<< metal4 >>
rect 565 885 595 1300
<< metal3 >>
rect 1310 1375 1354 1419
<< metal4 >>
rect 1310 1375 1354 1419
<< via3 >>
rect 1317 1382 1347 1412
<< metal3 >>
rect 1310 1263 1354 1307
<< metal4 >>
rect 1310 1263 1354 1307
<< via3 >>
rect 1317 1270 1347 1300
<< metal3 >>
rect 1902 1263 1946 1307
<< metal4 >>
rect 1902 1263 1946 1307
<< via3 >>
rect 1909 1270 1939 1300
<< metal3 >>
rect 1902 2063 1946 2107
<< metal4 >>
rect 1902 2063 1946 2107
<< via3 >>
rect 1909 2070 1939 2100
<< metal3 >>
rect 1310 2063 1354 2107
<< metal4 >>
rect 1310 2063 1354 2107
<< via3 >>
rect 1317 2070 1347 2100
<< metal3 >>
rect 1310 2559 1354 2603
<< metal4 >>
rect 1310 2559 1354 2603
<< via3 >>
rect 1317 2566 1347 2596
<< metal3 >>
rect 558 2559 602 2603
<< metal4 >>
rect 558 2559 602 2603
<< via3 >>
rect 565 2566 595 2596
<< metal3 >>
rect 558 2063 602 2107
<< metal4 >>
rect 558 2063 602 2107
<< via3 >>
rect 565 2070 595 2100
<< metal3 >>
rect 206 2063 250 2107
<< metal4 >>
rect 206 2063 250 2107
<< via3 >>
rect 213 2070 243 2100
<< metal3 >>
rect 206 1263 250 1307
<< metal4 >>
rect 206 1263 250 1307
<< via3 >>
rect 213 1270 243 1300
<< metal3 >>
rect 558 1263 602 1307
<< metal4 >>
rect 558 1263 602 1307
<< via3 >>
rect 565 1270 595 1300
<< metal4 >>
rect 5254 937 5284 1576
<< metal3 >>
rect 1190 1546 5284 1576
<< metal3 >>
rect 453 1546 1220 1576
<< metal3 >>
rect 5247 1539 5291 1583
<< metal4 >>
rect 5247 1539 5291 1583
<< via3 >>
rect 5254 1546 5284 1576
<< metal3 >>
rect 2243 921 4962 951
<< metal4 >>
rect 4932 921 4962 2807
<< metal3 >>
rect 4932 2777 5267 2807
<< metal3 >>
rect 4925 914 4969 958
<< metal4 >>
rect 4925 914 4969 958
<< via3 >>
rect 4932 921 4962 951
<< metal3 >>
rect 4925 2770 4969 2814
<< metal4 >>
rect 4925 2770 4969 2814
<< via3 >>
rect 4932 2777 4962 2807
<< metal4 >>
rect 2228 2011 2258 2794
<< metal3 >>
rect 2228 2011 5282 2041
<< metal4 >>
rect 5252 1866 5282 2041
<< metal3 >>
rect 2221 2004 2265 2048
<< metal4 >>
rect 2221 2004 2265 2048
<< via3 >>
rect 2228 2011 2258 2041
<< metal3 >>
rect 5245 2004 5289 2048
<< metal4 >>
rect 5245 2004 5289 2048
<< via3 >>
rect 5252 2011 5282 2041
<< metal1 >>
rect 100 3730 5586 3780
<< metal1 >>
rect 100 100 5586 150
<< metal2 >>
rect 100 150 150 3730
<< metal2 >>
rect 5536 150 5586 3730
<< metal1 >>
rect 93 3723 157 3787
<< metal2 >>
rect 93 3723 157 3787
<< via1 >>
rect 100 3730 150 3780
<< metal1 >>
rect 93 93 157 157
<< metal2 >>
rect 93 93 157 157
<< via1 >>
rect 100 100 150 150
<< metal1 >>
rect 5529 3723 5593 3787
<< metal2 >>
rect 5529 3723 5593 3787
<< via1 >>
rect 5536 3730 5586 3780
<< metal1 >>
rect 5529 93 5593 157
<< metal2 >>
rect 5529 93 5593 157
<< via1 >>
rect 5536 100 5586 150
<< metal1 >>
rect 0 3830 5686 3880
<< metal1 >>
rect 0 0 5686 50
<< metal2 >>
rect 0 50 50 3830
<< metal2 >>
rect 5636 50 5686 3830
<< metal1 >>
rect -7 3823 57 3887
<< metal2 >>
rect -7 3823 57 3887
<< via1 >>
rect 0 3830 50 3880
<< metal1 >>
rect -7 -7 57 57
<< metal2 >>
rect -7 -7 57 57
<< via1 >>
rect 0 0 50 50
<< metal1 >>
rect 5629 3823 5693 3887
<< metal2 >>
rect 5629 3823 5693 3887
<< via1 >>
rect 5636 3830 5686 3880
<< metal1 >>
rect 5629 -7 5693 57
<< metal2 >>
rect 5629 -7 5693 57
<< via1 >>
rect 5636 0 5686 50
<< metal1 >>
rect 2046 1850 2343 1890
<< metal1 >>
rect 2038 1024 5586 1080
<< metal1 >>
rect 5529 1017 5593 1087
<< metal2 >>
rect 5529 1017 5593 1087
<< via1 >>
rect 5536 1024 5586 1080
<< metal1 >>
rect 2038 200 5586 256
<< metal1 >>
rect 5529 193 5593 263
<< metal2 >>
rect 5529 193 5593 263
<< via1 >>
rect 5536 200 5586 256
<< metal1 >>
rect 2038 2884 5586 2940
<< metal1 >>
rect 5529 2877 5593 2947
<< metal2 >>
rect 5529 2877 5593 2947
<< via1 >>
rect 5536 2884 5586 2940
<< metal1 >>
rect 2038 2060 5586 2116
<< metal1 >>
rect 5529 2053 5593 2123
<< metal2 >>
rect 5529 2053 5593 2123
<< via1 >>
rect 5536 2060 5586 2116
<< metal1 >>
rect 2038 1954 5586 2010
<< metal1 >>
rect 5529 1947 5593 2017
<< metal2 >>
rect 5529 1947 5593 2017
<< via1 >>
rect 5536 1954 5586 2010
<< metal1 >>
rect 2038 1130 5586 1186
<< metal1 >>
rect 5529 1123 5593 1193
<< metal2 >>
rect 5529 1123 5593 1193
<< via1 >>
rect 5536 1130 5586 1186
<< metal1 >>
rect 1019 1664 1397 1704
<< metal1 >>
rect 263 1664 641 1704
<< metal1 >>
rect 767 1544 977 1584
<< metal1 >>
rect 1019 3580 1397 3620
<< metal1 >>
rect 1523 3460 1733 3500
<< metal1 >>
rect 263 3580 641 3620
<< metal1 >>
rect 0 2221 2132 2347
<< metal1 >>
rect -7 2214 57 2354
<< metal2 >>
rect -7 2214 57 2354
<< via1 >>
rect 0 2221 50 2347
<< metal1 >>
rect 0 2721 2132 2847
<< metal1 >>
rect -7 2714 57 2854
<< metal2 >>
rect -7 2714 57 2854
<< via1 >>
rect 0 2721 50 2847
<< metal1 >>
rect 0 2081 2132 2207
<< metal1 >>
rect -7 2074 57 2214
<< metal2 >>
rect -7 2074 57 2214
<< via1 >>
rect 0 2081 50 2207
<< metal1 >>
rect 0 381 2132 507
<< metal1 >>
rect -7 374 57 514
<< metal2 >>
rect -7 374 57 514
<< via1 >>
rect 0 381 50 507
<< metal1 >>
rect 100 3737 1964 3863
<< metal1 >>
rect 93 3730 157 3870
<< metal2 >>
rect 93 3730 157 3870
<< via1 >>
rect 100 3737 150 3863
<< metal1 >>
rect 100 3097 1964 3223
<< metal1 >>
rect 93 3090 157 3230
<< metal2 >>
rect 93 3090 157 3230
<< via1 >>
rect 100 3097 150 3223
<< metal2 >>
rect 424 1137 480 1191
<< metal3 >>
rect 424 1137 480 1191
<< via2 >>
rect 431 1144 473 1184
<< metal2 >>
rect 1180 1137 1236 1191
<< metal3 >>
rect 1180 1137 1236 1191
<< via2 >>
rect 1187 1144 1229 1184
<< metal2 >>
rect 1180 1137 1236 1191
<< metal3 >>
rect 1180 1137 1236 1191
<< via2 >>
rect 1187 1144 1229 1184
<< metal2 >>
rect 1180 1937 1236 1991
<< metal3 >>
rect 1180 1937 1236 1991
<< via2 >>
rect 1187 1944 1229 1984
<< metal2 >>
rect 1180 1937 1236 1991
<< metal3 >>
rect 1180 1937 1236 1991
<< via2 >>
rect 1187 1944 1229 1984
<< metal2 >>
rect 424 1937 480 1991
<< metal3 >>
rect 424 1937 480 1991
<< via2 >>
rect 431 1944 473 1984
<< metal2 >>
rect 1180 2437 1236 2491
<< metal3 >>
rect 1180 2437 1236 2491
<< via2 >>
rect 1187 2444 1229 2484
<< metal2 >>
rect 424 2437 480 2491
<< metal3 >>
rect 424 2437 480 2491
<< via2 >>
rect 431 2444 473 2484
<< metal2 >>
rect 424 2437 480 2491
<< metal3 >>
rect 424 2437 480 2491
<< via2 >>
rect 431 2444 473 2484
<< metal2 >>
rect 1180 737 1236 791
<< metal3 >>
rect 1180 737 1236 791
<< via2 >>
rect 1187 744 1229 784
<< metal2 >>
rect 424 737 480 791
<< metal3 >>
rect 424 737 480 791
<< via2 >>
rect 431 744 473 784
<< metal2 >>
rect 424 737 480 791
<< metal3 >>
rect 424 737 480 791
<< via2 >>
rect 431 744 473 784
<< metal2 >>
rect 1516 2277 1656 2331
<< metal3 >>
rect 1516 2277 1656 2331
<< via2 >>
rect 1523 2284 1649 2324
<< metal2 >>
rect 1516 2277 1656 2331
<< metal3 >>
rect 1516 2277 1656 2331
<< via2 >>
rect 1523 2284 1649 2324
<< metal2 >>
rect 760 2277 900 2331
<< metal3 >>
rect 760 2277 900 2331
<< metal4 >>
rect 760 2277 900 2331
<< via3 >>
rect 767 2284 893 2324
<< via2 >>
rect 767 2284 893 2324
<< metal2 >>
rect 760 2277 900 2331
<< metal3 >>
rect 760 2277 900 2331
<< via2 >>
rect 767 2284 893 2324
<< metal2 >>
rect 1516 577 1656 631
<< metal3 >>
rect 1516 577 1656 631
<< via2 >>
rect 1523 584 1649 624
<< metal2 >>
rect 1516 577 1656 631
<< metal3 >>
rect 1516 577 1656 631
<< via2 >>
rect 1523 584 1649 624
<< metal2 >>
rect 760 577 900 631
<< metal3 >>
rect 760 577 900 631
<< via2 >>
rect 767 584 893 624
<< metal2 >>
rect 760 3293 900 3347
<< metal3 >>
rect 760 3293 900 3347
<< metal4 >>
rect 760 3293 900 3347
<< via3 >>
rect 767 3300 893 3340
<< via2 >>
rect 767 3300 893 3340
<< metal2 >>
rect 760 977 900 1031
<< metal3 >>
rect 760 977 900 1031
<< via2 >>
rect 767 984 893 1024
<< metal2 >>
rect 1516 977 1656 1031
<< metal3 >>
rect 1516 977 1656 1031
<< via2 >>
rect 1523 984 1649 1024
<< metal2 >>
rect 1516 977 1656 1031
<< metal3 >>
rect 1516 977 1656 1031
<< via2 >>
rect 1523 984 1649 1024
<< metal2 >>
rect 1516 1777 1656 1831
<< metal3 >>
rect 1516 1777 1656 1831
<< via2 >>
rect 1523 1784 1649 1824
<< metal2 >>
rect 1516 1777 1656 1831
<< metal3 >>
rect 1516 1777 1656 1831
<< via2 >>
rect 1523 1784 1649 1824
<< metal2 >>
rect 760 1777 900 1831
<< metal3 >>
rect 760 1777 900 1831
<< via2 >>
rect 767 1784 893 1824
<< metal2 >>
rect 760 1777 900 1831
<< metal3 >>
rect 760 1777 900 1831
<< via2 >>
rect 767 1784 893 1824
<< metal2 >>
rect 1180 3453 1236 3507
<< metal3 >>
rect 1180 3453 1236 3507
<< via2 >>
rect 1187 3460 1229 3500
<< metal2 >>
rect 424 3453 480 3507
<< metal3 >>
rect 424 3453 480 3507
<< via2 >>
rect 431 3460 473 3500
<< metal2 >>
rect 424 3453 480 3507
<< metal3 >>
rect 424 3453 480 3507
<< via2 >>
rect 431 3460 473 3500
<< metal2 >>
rect 508 1257 648 1311
<< metal3 >>
rect 508 1257 648 1311
<< via2 >>
rect 515 1264 641 1304
<< metal2 >>
rect 508 1257 648 1311
<< metal3 >>
rect 508 1257 648 1311
<< metal4 >>
rect 508 1257 648 1311
<< via3 >>
rect 515 1264 641 1304
<< via2 >>
rect 515 1264 641 1304
<< metal2 >>
rect 1264 1257 1404 1311
<< metal3 >>
rect 1264 1257 1404 1311
<< metal4 >>
rect 1264 1257 1404 1311
<< via3 >>
rect 1271 1264 1397 1304
<< via2 >>
rect 1271 1264 1397 1304
<< metal2 >>
rect 1264 1257 1404 1311
<< metal3 >>
rect 1264 1257 1404 1311
<< metal4 >>
rect 1264 1257 1404 1311
<< via3 >>
rect 1271 1264 1397 1304
<< via2 >>
rect 1271 1264 1397 1304
<< metal2 >>
rect 1264 1257 1404 1311
<< metal3 >>
rect 1264 1257 1404 1311
<< via2 >>
rect 1271 1264 1397 1304
<< metal2 >>
rect 1264 2057 1404 2111
<< metal3 >>
rect 1264 2057 1404 2111
<< via2 >>
rect 1271 2064 1397 2104
<< metal2 >>
rect 1264 2057 1404 2111
<< metal3 >>
rect 1264 2057 1404 2111
<< metal4 >>
rect 1264 2057 1404 2111
<< via3 >>
rect 1271 2064 1397 2104
<< via2 >>
rect 1271 2064 1397 2104
<< metal2 >>
rect 508 2057 648 2111
<< metal3 >>
rect 508 2057 648 2111
<< metal4 >>
rect 508 2057 648 2111
<< via3 >>
rect 515 2064 641 2104
<< via2 >>
rect 515 2064 641 2104
<< metal2 >>
rect 508 2057 648 2111
<< metal3 >>
rect 508 2057 648 2111
<< via2 >>
rect 515 2064 641 2104
<< metal2 >>
rect 1264 2557 1404 2611
<< metal3 >>
rect 1264 2557 1404 2611
<< metal4 >>
rect 1264 2557 1404 2611
<< via3 >>
rect 1271 2564 1397 2604
<< via2 >>
rect 1271 2564 1397 2604
<< metal2 >>
rect 1264 2557 1404 2611
<< metal3 >>
rect 1264 2557 1404 2611
<< via2 >>
rect 1271 2564 1397 2604
<< metal2 >>
rect 508 2557 648 2611
<< metal3 >>
rect 508 2557 648 2611
<< via2 >>
rect 515 2564 641 2604
<< metal2 >>
rect 508 2557 648 2611
<< metal3 >>
rect 508 2557 648 2611
<< metal4 >>
rect 508 2557 648 2611
<< via3 >>
rect 515 2564 641 2604
<< via2 >>
rect 515 2564 641 2604
<< metal2 >>
rect 1264 857 1404 911
<< metal3 >>
rect 1264 857 1404 911
<< metal4 >>
rect 1264 857 1404 911
<< via3 >>
rect 1271 864 1397 904
<< via2 >>
rect 1271 864 1397 904
<< metal2 >>
rect 1264 857 1404 911
<< metal3 >>
rect 1264 857 1404 911
<< metal4 >>
rect 1264 857 1404 911
<< via3 >>
rect 1271 864 1397 904
<< via2 >>
rect 1271 864 1397 904
<< metal2 >>
rect 508 857 648 911
<< metal3 >>
rect 508 857 648 911
<< metal4 >>
rect 508 857 648 911
<< via3 >>
rect 515 864 641 904
<< via2 >>
rect 515 864 641 904
<< metal2 >>
rect 1516 1377 1656 1431
<< metal3 >>
rect 1516 1377 1656 1431
<< via2 >>
rect 1523 1384 1649 1424
<< metal2 >>
rect 1180 1537 1236 1591
<< metal3 >>
rect 1180 1537 1236 1591
<< via2 >>
rect 1187 1544 1229 1584
<< metal2 >>
rect 1180 1537 1236 1591
<< metal3 >>
rect 1180 1537 1236 1591
<< via2 >>
rect 1187 1544 1229 1584
<< metal2 >>
rect 424 1537 480 1591
<< metal3 >>
rect 424 1537 480 1591
<< via2 >>
rect 431 1544 473 1584
<< metal1 >>
rect 5174 913 5386 967
<< metal2 >>
rect 5174 913 5386 967
<< metal3 >>
rect 5174 913 5386 967
<< metal4 >>
rect 5174 913 5386 967
<< via3 >>
rect 5181 920 5379 960
<< via2 >>
rect 5181 920 5379 960
<< via1 >>
rect 5181 920 5379 960
<< metal1 >>
rect 2138 913 2350 967
<< metal2 >>
rect 2138 913 2350 967
<< metal3 >>
rect 2138 913 2350 967
<< via2 >>
rect 2145 920 2343 960
<< via1 >>
rect 2145 920 2343 960
<< metal1 >>
rect 5174 2773 5386 2827
<< metal2 >>
rect 5174 2773 5386 2827
<< metal3 >>
rect 5174 2773 5386 2827
<< via2 >>
rect 5181 2780 5379 2820
<< via1 >>
rect 5181 2780 5379 2820
<< metal1 >>
rect 2138 2773 2350 2827
<< metal2 >>
rect 2138 2773 2350 2827
<< metal3 >>
rect 2138 2773 2350 2827
<< metal4 >>
rect 2138 2773 2350 2827
<< via3 >>
rect 2145 2780 2343 2820
<< via2 >>
rect 2145 2780 2343 2820
<< via1 >>
rect 2145 2780 2343 2820
<< metal1 >>
rect 5174 1843 5386 1897
<< metal2 >>
rect 5174 1843 5386 1897
<< metal3 >>
rect 5174 1843 5386 1897
<< metal4 >>
rect 5174 1843 5386 1897
<< via3 >>
rect 5181 1850 5379 1890
<< via2 >>
rect 5181 1850 5379 1890
<< via1 >>
rect 5181 1850 5379 1890
<< labels >>
flabel metal3 s 454 1947 1221 1977 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel metal3 s 439 749 1206 779 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel metal1 s 0 3830 5686 3880 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel metal1 s 100 3730 5586 3780 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel metal4 s 808 2285 838 3324 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>