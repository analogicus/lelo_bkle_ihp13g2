magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747405728
<< checkpaint >>
rect 0 0 1 1
use LELOTR_NCHDL  None_MN2 ../LELO_TR_IHP13G2
timestamp 1747405728
transform 1 0 200 0 1 200
box 0 0 407 160
use LELOTR_NCHDL  None_MN3 ../LELO_TR_IHP13G2
timestamp 1747405728
transform 1 0 607 0 1 200
box 0 0 407 160
use LELOTR_PCHDL  None_MP2 ../LELO_TR_IHP13G2
timestamp 1747405728
transform 1 0 607 0 1 1080
box 0 0 407 160
use LELOTR_PCHDL  None_MP3 ../LELO_TR_IHP13G2
timestamp 1747405728
transform 1 0 200 0 1 1080
box 0 0 407 160
<< metal4 >>
rect 327 278 357 1029
<< metal3 >>
rect 327 999 885 1029
<< metal4 >>
rect 855 999 885 1158
<< metal3 >>
rect 320 992 364 1036
<< metal4 >>
rect 320 992 364 1036
<< via3 >>
rect 327 999 357 1029
<< metal3 >>
rect 848 992 892 1036
<< metal4 >>
rect 848 992 892 1036
<< via3 >>
rect 855 999 885 1029
<< metal4 >>
rect 730 278 760 917
<< metal3 >>
rect 442 887 760 917
<< metal4 >>
rect 442 887 472 1158
<< metal3 >>
rect 723 880 767 924
<< metal4 >>
rect 723 880 767 924
<< via3 >>
rect 730 887 760 917
<< metal3 >>
rect 435 880 479 924
<< metal4 >>
rect 435 880 479 924
<< via3 >>
rect 442 887 472 917
<< metal3 >>
rect 169 1101 312 1131
<< metal4 >>
rect 169 429 199 1131
<< metal3 >>
rect 169 429 919 459
<< metal4 >>
rect 889 301 919 459
<< metal4 >>
rect 889 301 919 795
<< metal3 >>
rect 569 765 919 795
<< metal4 >>
rect 569 765 599 1211
<< metal3 >>
rect 569 1181 712 1211
<< metal3 >>
rect 162 1094 206 1138
<< metal4 >>
rect 162 1094 206 1138
<< via3 >>
rect 169 1101 199 1131
<< metal3 >>
rect 162 422 206 466
<< metal4 >>
rect 162 422 206 466
<< via3 >>
rect 169 429 199 459
<< metal3 >>
rect 882 422 926 466
<< metal4 >>
rect 882 422 926 466
<< via3 >>
rect 889 429 919 459
<< metal3 >>
rect 882 758 926 802
<< metal4 >>
rect 882 758 926 802
<< via3 >>
rect 889 765 919 795
<< metal3 >>
rect 562 758 606 802
<< metal4 >>
rect 562 758 606 802
<< via3 >>
rect 569 765 599 795
<< metal3 >>
rect 562 1174 606 1218
<< metal4 >>
rect 562 1174 606 1218
<< via3 >>
rect 569 1181 599 1211
<< metal1 >>
rect 100 1290 1114 1340
<< metal1 >>
rect 100 100 1114 150
<< metal2 >>
rect 100 150 150 1290
<< metal2 >>
rect 1064 150 1114 1290
<< metal1 >>
rect 93 1283 157 1347
<< metal2 >>
rect 93 1283 157 1347
<< via1 >>
rect 100 1290 150 1340
<< metal1 >>
rect 93 93 157 157
<< metal2 >>
rect 93 93 157 157
<< via1 >>
rect 100 100 150 150
<< metal1 >>
rect 1057 1283 1121 1347
<< metal2 >>
rect 1057 1283 1121 1347
<< via1 >>
rect 1064 1290 1114 1340
<< metal1 >>
rect 1057 93 1121 157
<< metal2 >>
rect 1057 93 1121 157
<< via1 >>
rect 1064 100 1114 150
<< metal1 >>
rect 0 1390 1214 1440
<< metal1 >>
rect 0 0 1214 50
<< metal2 >>
rect 0 50 50 1390
<< metal2 >>
rect 1164 50 1214 1390
<< metal1 >>
rect -7 1383 57 1447
<< metal2 >>
rect -7 1383 57 1447
<< via1 >>
rect 0 1390 50 1440
<< metal1 >>
rect -7 -7 57 57
<< metal2 >>
rect -7 -7 57 57
<< via1 >>
rect 0 0 50 50
<< metal1 >>
rect 1157 1383 1221 1447
<< metal2 >>
rect 1157 1383 1221 1447
<< via1 >>
rect 1164 1390 1214 1440
<< metal1 >>
rect 1157 -7 1221 57
<< metal2 >>
rect 1157 -7 1221 57
<< via1 >>
rect 1164 0 1214 50
<< metal1 >>
rect 292 263 394 297
<< metal2 >>
rect 292 263 394 297
<< metal3 >>
rect 292 263 394 297
<< metal4 >>
rect 292 263 394 297
<< via3 >>
rect 299 270 387 290
<< via2 >>
rect 299 270 387 290
<< via1 >>
rect 299 270 387 290
<< metal1 >>
rect 820 1143 922 1177
<< metal2 >>
rect 820 1143 922 1177
<< metal3 >>
rect 820 1143 922 1177
<< metal4 >>
rect 820 1143 922 1177
<< via3 >>
rect 827 1150 915 1170
<< via2 >>
rect 827 1150 915 1170
<< via1 >>
rect 827 1150 915 1170
<< metal1 >>
rect 699 263 801 297
<< metal2 >>
rect 699 263 801 297
<< metal3 >>
rect 699 263 801 297
<< metal4 >>
rect 699 263 801 297
<< via3 >>
rect 706 270 794 290
<< via2 >>
rect 706 270 794 290
<< via1 >>
rect 706 270 794 290
<< metal1 >>
rect 413 1143 515 1177
<< metal2 >>
rect 413 1143 515 1177
<< metal3 >>
rect 413 1143 515 1177
<< metal4 >>
rect 413 1143 515 1177
<< via3 >>
rect 420 1150 508 1170
<< via2 >>
rect 420 1150 508 1170
<< via1 >>
rect 420 1150 508 1170
<< metal1 >>
rect 853 303 955 337
<< metal2 >>
rect 853 303 955 337
<< metal3 >>
rect 853 303 955 337
<< metal4 >>
rect 853 303 955 337
<< via3 >>
rect 860 310 948 330
<< via2 >>
rect 860 310 948 330
<< via1 >>
rect 860 310 948 330
<< metal1 >>
rect 853 303 955 337
<< metal2 >>
rect 853 303 955 337
<< metal3 >>
rect 853 303 955 337
<< metal4 >>
rect 853 303 955 337
<< via3 >>
rect 860 310 948 330
<< via2 >>
rect 860 310 948 330
<< via1 >>
rect 860 310 948 330
<< metal1 >>
rect 666 1183 768 1217
<< metal2 >>
rect 666 1183 768 1217
<< metal3 >>
rect 666 1183 768 1217
<< via2 >>
rect 673 1190 761 1210
<< via1 >>
rect 673 1190 761 1210
<< metal1 >>
rect 259 1103 361 1137
<< metal2 >>
rect 259 1103 361 1137
<< metal3 >>
rect 259 1103 361 1137
<< via2 >>
rect 266 1110 354 1130
<< via1 >>
rect 266 1110 354 1130
<< labels >>
flabel metal4 s 327 278 357 1029 0 FreeSans 400 0 0 0 A
port 23 nsew signal bidirectional
flabel metal4 s 730 278 760 917 0 FreeSans 400 0 0 0 B
port 24 nsew signal bidirectional
flabel metal3 s 169 1101 312 1131 0 FreeSans 400 0 0 0 Y
port 25 nsew signal bidirectional
flabel metal1 s 0 1390 1214 1440 0 FreeSans 400 0 0 0 AVDD
port 26 nsew signal bidirectional
flabel metal1 s 100 1290 1114 1340 0 FreeSans 400 0 0 0 AVSS
port 27 nsew signal bidirectional
<< properties >>
<< end >>