magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747934190
<< checkpaint >>
rect 0 0 1 1
use LELOATR_PCH_4C5F0  diff1_MP3<3> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 1450
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP3<2> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 1450
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP3<1> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 1850
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP3<0> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 1850
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP4<3> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 650
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  diff1_MP4<3>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 410
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<2> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 650
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  diff1_MP4<2>_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 410
box 0 0 756 240
use LELOATR_PCH_4C5F0  diff1_MP4<1> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 1050
box 0 0 756 400
use LELOATR_PCH_4C5F0  diff1_MP4<0> ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 1050
box 0 0 756 400
use LELOATR_PCH_4C5F0  mirror1_MP2 ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 2250
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  mirror1_MP2_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 2650
box 0 0 756 240
use LELOATR_PCH_4C5F0  mirror1_MP1 ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 2250
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  mirror1_MP1_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 2650
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN1 ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 3266
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN1_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 3666
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror2_MN1_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 3808 0 1 3026
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN2 ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 3266
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN2_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 3666
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror2_MN2_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747934190
transform 1 0 4564 0 1 3026
box 0 0 756 240
use LELOTR_RPPO16  bias1_RH1 ../LELO_TR_IHP13G2
timestamp 1747934190
transform 1 0 160 0 1 200
box 0 0 3448 880
use LELOTR_RPPO16  bias1_RH2 ../LELO_TR_IHP13G2
timestamp 1747934190
transform 1 0 160 0 1 2060
box 0 0 3448 880
use LELOTR_RPPO16  bias1_RH3 ../LELO_TR_IHP13G2
timestamp 1747934190
transform 1 0 160 0 1 1130
box 0 0 3448 880
<< metal3 >>
rect 4543 1631 4686 1661
<< metal4 >>
rect 4543 1631 4573 2061
<< metal3 >>
rect 4543 2031 4701 2061
<< metal3 >>
rect 3919 2031 4701 2061
<< metal3 >>
rect 3791 2031 3949 2061
<< metal4 >>
rect 3791 1631 3821 2061
<< metal3 >>
rect 3791 1631 3934 1661
<< metal3 >>
rect 4536 1624 4580 1668
<< metal4 >>
rect 4536 1624 4580 1668
<< via3 >>
rect 4543 1631 4573 1661
<< metal3 >>
rect 4536 2024 4580 2068
<< metal4 >>
rect 4536 2024 4580 2068
<< via3 >>
rect 4543 2031 4573 2061
<< metal3 >>
rect 3784 2024 3828 2068
<< metal4 >>
rect 3784 2024 3828 2068
<< via3 >>
rect 3791 2031 3821 2061
<< metal3 >>
rect 3784 1624 3828 1668
<< metal4 >>
rect 3784 1624 3828 1668
<< via3 >>
rect 3791 1631 3821 1661
<< metal3 >>
rect 3791 831 3934 861
<< metal4 >>
rect 3791 831 3821 1261
<< metal3 >>
rect 3791 1231 3949 1261
<< metal3 >>
rect 3919 1231 4701 1261
<< metal3 >>
rect 4543 1231 4701 1261
<< metal4 >>
rect 4543 831 4573 1261
<< metal3 >>
rect 4543 831 4686 861
<< metal3 >>
rect 3784 824 3828 868
<< metal4 >>
rect 3784 824 3828 868
<< via3 >>
rect 3791 831 3821 861
<< metal3 >>
rect 3784 1224 3828 1268
<< metal4 >>
rect 3784 1224 3828 1268
<< via3 >>
rect 3791 1231 3821 1261
<< metal3 >>
rect 4536 1224 4580 1268
<< metal4 >>
rect 4536 1224 4580 1268
<< via3 >>
rect 4543 1231 4573 1261
<< metal3 >>
rect 4536 824 4580 868
<< metal4 >>
rect 4536 824 4580 868
<< via3 >>
rect 4543 831 4573 861
<< metal3 >>
rect 5073 3296 5232 3326
<< metal4 >>
rect 5202 1072 5232 3326
<< metal3 >>
rect 5058 1072 5232 1102
<< metal4 >>
rect 5058 672 5088 1102
<< metal3 >>
rect 4290 672 5088 702
<< metal4 >>
rect 4290 672 4320 1087
<< metal3 >>
rect 5195 3289 5239 3333
<< metal4 >>
rect 5195 3289 5239 3333
<< via3 >>
rect 5202 3296 5232 3326
<< metal3 >>
rect 5195 1065 5239 1109
<< metal4 >>
rect 5195 1065 5239 1109
<< via3 >>
rect 5202 1072 5232 1102
<< metal3 >>
rect 5051 1065 5095 1109
<< metal4 >>
rect 5051 1065 5095 1109
<< via3 >>
rect 5058 1072 5088 1102
<< metal3 >>
rect 5051 665 5095 709
<< metal4 >>
rect 5051 665 5095 709
<< via3 >>
rect 5058 672 5088 702
<< metal3 >>
rect 4283 665 4327 709
<< metal4 >>
rect 4283 665 4327 709
<< via3 >>
rect 4290 672 4320 702
<< metal3 >>
rect 3921 3455 4688 3485
<< metal3 >>
rect 3921 3455 4463 3485
<< metal4 >>
rect 4433 1871 4463 3485
<< metal3 >>
rect 4289 1871 4463 1901
<< metal4 >>
rect 4289 1471 4319 1901
<< metal3 >>
rect 4289 1471 5087 1501
<< metal4 >>
rect 5057 1471 5087 1886
<< metal3 >>
rect 4426 3448 4470 3492
<< metal4 >>
rect 4426 3448 4470 3492
<< via3 >>
rect 4433 3455 4463 3485
<< metal3 >>
rect 4426 1864 4470 1908
<< metal4 >>
rect 4426 1864 4470 1908
<< via3 >>
rect 4433 1871 4463 1901
<< metal3 >>
rect 4282 1864 4326 1908
<< metal4 >>
rect 4282 1864 4326 1908
<< via3 >>
rect 4289 1871 4319 1901
<< metal3 >>
rect 4282 1464 4326 1508
<< metal4 >>
rect 4282 1464 4326 1508
<< via3 >>
rect 4289 1471 4319 1501
<< metal3 >>
rect 5050 1464 5094 1508
<< metal4 >>
rect 5050 1464 5094 1508
<< via3 >>
rect 5057 1471 5087 1501
<< metal3 >>
rect 4799 2266 5070 2296
<< metal4 >>
rect 4799 1769 4829 2296
<< metal3 >>
rect 4792 2259 4836 2303
<< metal4 >>
rect 4792 2259 4836 2303
<< via3 >>
rect 4799 2266 4829 2296
<< metal3 >>
rect 3391 926 3678 956
<< metal4 >>
rect 3648 926 3678 2460
<< metal3 >>
rect 3648 2430 3950 2460
<< metal3 >>
rect 3920 2430 4687 2460
<< metal3 >>
rect 3641 919 3685 963
<< metal4 >>
rect 3641 919 3685 963
<< via3 >>
rect 3648 926 3678 956
<< metal3 >>
rect 3641 2423 3685 2467
<< metal4 >>
rect 3641 2423 3685 2467
<< via3 >>
rect 3648 2430 3678 2460
<< metal3 >>
rect 365 921 3164 951
<< metal4 >>
rect 3134 921 3164 2807
<< metal3 >>
rect 3134 2777 3389 2807
<< metal3 >>
rect 3127 914 3171 958
<< metal4 >>
rect 3127 914 3171 958
<< via3 >>
rect 3134 921 3164 951
<< metal3 >>
rect 3127 2770 3171 2814
<< metal4 >>
rect 3127 2770 3171 2814
<< via3 >>
rect 3134 2777 3164 2807
<< metal4 >>
rect 350 1995 380 2794
<< metal3 >>
rect 350 1995 3404 2025
<< metal4 >>
rect 3374 1866 3404 2025
<< metal3 >>
rect 343 1988 387 2032
<< metal4 >>
rect 343 1988 387 2032
<< via3 >>
rect 350 1995 380 2025
<< metal3 >>
rect 3367 1988 3411 2032
<< metal4 >>
rect 3367 1988 3411 2032
<< via3 >>
rect 3374 1995 3404 2025
<< metal1 >>
rect 100 3956 5500 4006
<< metal1 >>
rect 100 100 5500 150
<< metal2 >>
rect 100 150 150 3956
<< metal2 >>
rect 5450 150 5500 3956
<< metal1 >>
rect 93 3949 157 4013
<< metal2 >>
rect 93 3949 157 4013
<< via1 >>
rect 100 3956 150 4006
<< metal1 >>
rect 93 93 157 157
<< metal2 >>
rect 93 93 157 157
<< via1 >>
rect 100 100 150 150
<< metal1 >>
rect 5443 3949 5507 4013
<< metal2 >>
rect 5443 3949 5507 4013
<< via1 >>
rect 5450 3956 5500 4006
<< metal1 >>
rect 5443 93 5507 157
<< metal2 >>
rect 5443 93 5507 157
<< via1 >>
rect 5450 100 5500 150
<< metal1 >>
rect 0 4056 5600 4106
<< metal1 >>
rect 0 0 5600 50
<< metal2 >>
rect 0 50 50 4056
<< metal2 >>
rect 5550 50 5600 4056
<< metal1 >>
rect -7 4049 57 4113
<< metal2 >>
rect -7 4049 57 4113
<< via1 >>
rect 0 4056 50 4106
<< metal1 >>
rect -7 -7 57 57
<< metal2 >>
rect -7 -7 57 57
<< via1 >>
rect 0 0 50 50
<< metal1 >>
rect 5543 4049 5607 4113
<< metal2 >>
rect 5543 4049 5607 4113
<< via1 >>
rect 5550 4056 5600 4106
<< metal1 >>
rect 5543 -7 5607 57
<< metal2 >>
rect 5543 -7 5607 57
<< via1 >>
rect 5550 0 5600 50
<< metal1 >>
rect 168 1850 465 1890
<< metal1 >>
rect 100 1024 3548 1080
<< metal1 >>
rect 93 1017 157 1087
<< metal2 >>
rect 93 1017 157 1087
<< via1 >>
rect 100 1024 150 1080
<< metal1 >>
rect 100 200 3548 256
<< metal1 >>
rect 93 193 157 263
<< metal2 >>
rect 93 193 157 263
<< via1 >>
rect 100 200 150 256
<< metal1 >>
rect 100 2884 3548 2940
<< metal1 >>
rect 93 2877 157 2947
<< metal2 >>
rect 93 2877 157 2947
<< via1 >>
rect 100 2884 150 2940
<< metal1 >>
rect 100 2060 3548 2116
<< metal1 >>
rect 93 2053 157 2123
<< metal2 >>
rect 93 2053 157 2123
<< via1 >>
rect 100 2060 150 2116
<< metal1 >>
rect 100 1954 3548 2010
<< metal1 >>
rect 93 1947 157 2017
<< metal2 >>
rect 93 1947 157 2017
<< via1 >>
rect 100 1954 150 2010
<< metal1 >>
rect 100 1130 3548 1186
<< metal1 >>
rect 93 1123 157 1193
<< metal2 >>
rect 93 1123 157 1193
<< via1 >>
rect 100 1130 150 1186
<< metal1 >>
rect 4501 2550 4879 2590
<< metal1 >>
rect 3745 2550 4123 2590
<< metal1 >>
rect 4249 2430 4459 2470
<< metal1 >>
rect 3745 3566 4123 3606
<< metal1 >>
rect 4249 3446 4459 3486
<< metal1 >>
rect 4501 3566 4879 3606
<< metal1 >>
rect 3888 467 5600 593
<< metal1 >>
rect 5543 460 5607 600
<< metal2 >>
rect 5543 460 5607 600
<< via1 >>
rect 5550 467 5600 593
<< metal1 >>
rect 3888 2707 5600 2833
<< metal1 >>
rect 5543 2700 5607 2840
<< metal2 >>
rect 5543 2700 5607 2840
<< via1 >>
rect 5550 2707 5600 2833
<< metal1 >>
rect 3888 3723 5500 3849
<< metal1 >>
rect 5443 3716 5507 3856
<< metal2 >>
rect 5443 3716 5507 3856
<< via1 >>
rect 5450 3723 5500 3849
<< metal1 >>
rect 3888 3083 5500 3209
<< metal1 >>
rect 5443 3076 5507 3216
<< metal2 >>
rect 5443 3076 5507 3216
<< via1 >>
rect 5450 3083 5500 3209
<< metal2 >>
rect 3906 1623 3962 1677
<< metal3 >>
rect 3906 1623 3962 1677
<< via2 >>
rect 3913 1630 3955 1670
<< metal2 >>
rect 4662 1623 4718 1677
<< metal3 >>
rect 4662 1623 4718 1677
<< via2 >>
rect 4669 1630 4711 1670
<< metal2 >>
rect 3906 2023 3962 2077
<< metal3 >>
rect 3906 2023 3962 2077
<< via2 >>
rect 3913 2030 3955 2070
<< metal2 >>
rect 3906 2023 3962 2077
<< metal3 >>
rect 3906 2023 3962 2077
<< via2 >>
rect 3913 2030 3955 2070
<< metal2 >>
rect 4662 2023 4718 2077
<< metal3 >>
rect 4662 2023 4718 2077
<< via2 >>
rect 4669 2030 4711 2070
<< metal2 >>
rect 4662 2023 4718 2077
<< metal3 >>
rect 4662 2023 4718 2077
<< via2 >>
rect 4669 2030 4711 2070
<< metal2 >>
rect 4662 823 4718 877
<< metal3 >>
rect 4662 823 4718 877
<< via2 >>
rect 4669 830 4711 870
<< metal2 >>
rect 3906 823 3962 877
<< metal3 >>
rect 3906 823 3962 877
<< via2 >>
rect 3913 830 3955 870
<< metal2 >>
rect 3906 1223 3962 1277
<< metal3 >>
rect 3906 1223 3962 1277
<< via2 >>
rect 3913 1230 3955 1270
<< metal2 >>
rect 3906 1223 3962 1277
<< metal3 >>
rect 3906 1223 3962 1277
<< via2 >>
rect 3913 1230 3955 1270
<< metal2 >>
rect 4662 1223 4718 1277
<< metal3 >>
rect 4662 1223 4718 1277
<< via2 >>
rect 4669 1230 4711 1270
<< metal2 >>
rect 4662 1223 4718 1277
<< metal3 >>
rect 4662 1223 4718 1277
<< via2 >>
rect 4669 1230 4711 1270
<< metal2 >>
rect 4998 663 5138 717
<< metal3 >>
rect 4998 663 5138 717
<< metal4 >>
rect 4998 663 5138 717
<< via3 >>
rect 5005 670 5131 710
<< via2 >>
rect 5005 670 5131 710
<< metal2 >>
rect 4998 663 5138 717
<< metal3 >>
rect 4998 663 5138 717
<< via2 >>
rect 5005 670 5131 710
<< metal2 >>
rect 4242 663 4382 717
<< metal3 >>
rect 4242 663 4382 717
<< via2 >>
rect 4249 670 4375 710
<< metal2 >>
rect 4242 663 4382 717
<< metal3 >>
rect 4242 663 4382 717
<< metal4 >>
rect 4242 663 4382 717
<< via3 >>
rect 4249 670 4375 710
<< via2 >>
rect 4249 670 4375 710
<< metal2 >>
rect 4242 1063 4382 1117
<< metal3 >>
rect 4242 1063 4382 1117
<< metal4 >>
rect 4242 1063 4382 1117
<< via3 >>
rect 4249 1070 4375 1110
<< via2 >>
rect 4249 1070 4375 1110
<< metal2 >>
rect 4998 1063 5138 1117
<< metal3 >>
rect 4998 1063 5138 1117
<< via2 >>
rect 5005 1070 5131 1110
<< metal2 >>
rect 4998 1063 5138 1117
<< metal3 >>
rect 4998 1063 5138 1117
<< metal4 >>
rect 4998 1063 5138 1117
<< via3 >>
rect 5005 1070 5131 1110
<< via2 >>
rect 5005 1070 5131 1110
<< metal2 >>
rect 4998 3279 5138 3333
<< metal3 >>
rect 4998 3279 5138 3333
<< via2 >>
rect 5005 3286 5131 3326
<< metal2 >>
rect 4242 1463 4382 1517
<< metal3 >>
rect 4242 1463 4382 1517
<< metal4 >>
rect 4242 1463 4382 1517
<< via3 >>
rect 4249 1470 4375 1510
<< via2 >>
rect 4249 1470 4375 1510
<< metal2 >>
rect 4242 1463 4382 1517
<< metal3 >>
rect 4242 1463 4382 1517
<< via2 >>
rect 4249 1470 4375 1510
<< metal2 >>
rect 4998 1463 5138 1517
<< metal3 >>
rect 4998 1463 5138 1517
<< via2 >>
rect 5005 1470 5131 1510
<< metal2 >>
rect 4998 1463 5138 1517
<< metal3 >>
rect 4998 1463 5138 1517
<< metal4 >>
rect 4998 1463 5138 1517
<< via3 >>
rect 5005 1470 5131 1510
<< via2 >>
rect 5005 1470 5131 1510
<< metal2 >>
rect 4242 1863 4382 1917
<< metal3 >>
rect 4242 1863 4382 1917
<< via2 >>
rect 4249 1870 4375 1910
<< metal2 >>
rect 4242 1863 4382 1917
<< metal3 >>
rect 4242 1863 4382 1917
<< metal4 >>
rect 4242 1863 4382 1917
<< via3 >>
rect 4249 1870 4375 1910
<< via2 >>
rect 4249 1870 4375 1910
<< metal2 >>
rect 4998 1863 5138 1917
<< metal3 >>
rect 4998 1863 5138 1917
<< metal4 >>
rect 4998 1863 5138 1917
<< via3 >>
rect 5005 1870 5131 1910
<< via2 >>
rect 5005 1870 5131 1910
<< metal2 >>
rect 3906 3439 3962 3493
<< metal3 >>
rect 3906 3439 3962 3493
<< via2 >>
rect 3913 3446 3955 3486
<< metal2 >>
rect 3906 3439 3962 3493
<< metal3 >>
rect 3906 3439 3962 3493
<< via2 >>
rect 3913 3446 3955 3486
<< metal2 >>
rect 4662 3439 4718 3493
<< metal3 >>
rect 4662 3439 4718 3493
<< via2 >>
rect 4669 3446 4711 3486
<< metal2 >>
rect 4746 1743 4886 1797
<< metal3 >>
rect 4746 1743 4886 1797
<< metal4 >>
rect 4746 1743 4886 1797
<< via3 >>
rect 4753 1750 4879 1790
<< via2 >>
rect 4753 1750 4879 1790
<< metal2 >>
rect 4746 2143 4886 2197
<< metal3 >>
rect 4746 2143 4886 2197
<< metal4 >>
rect 4746 2143 4886 2197
<< via3 >>
rect 4753 2150 4879 2190
<< via2 >>
rect 4753 2150 4879 2190
<< metal2 >>
rect 4998 2263 5138 2317
<< metal3 >>
rect 4998 2263 5138 2317
<< via2 >>
rect 5005 2270 5131 2310
<< metal2 >>
rect 4662 2423 4718 2477
<< metal3 >>
rect 4662 2423 4718 2477
<< via2 >>
rect 4669 2430 4711 2470
<< metal2 >>
rect 3906 2423 3962 2477
<< metal3 >>
rect 3906 2423 3962 2477
<< via2 >>
rect 3913 2430 3955 2470
<< metal2 >>
rect 3906 2423 3962 2477
<< metal3 >>
rect 3906 2423 3962 2477
<< via2 >>
rect 3913 2430 3955 2470
<< metal1 >>
rect 3296 913 3508 967
<< metal2 >>
rect 3296 913 3508 967
<< metal3 >>
rect 3296 913 3508 967
<< via2 >>
rect 3303 920 3501 960
<< via1 >>
rect 3303 920 3501 960
<< metal1 >>
rect 260 913 472 967
<< metal2 >>
rect 260 913 472 967
<< metal3 >>
rect 260 913 472 967
<< via2 >>
rect 267 920 465 960
<< via1 >>
rect 267 920 465 960
<< metal1 >>
rect 3296 2773 3508 2827
<< metal2 >>
rect 3296 2773 3508 2827
<< metal3 >>
rect 3296 2773 3508 2827
<< via2 >>
rect 3303 2780 3501 2820
<< via1 >>
rect 3303 2780 3501 2820
<< metal1 >>
rect 260 2773 472 2827
<< metal2 >>
rect 260 2773 472 2827
<< metal3 >>
rect 260 2773 472 2827
<< metal4 >>
rect 260 2773 472 2827
<< via3 >>
rect 267 2780 465 2820
<< via2 >>
rect 267 2780 465 2820
<< via1 >>
rect 267 2780 465 2820
<< metal1 >>
rect 3296 1843 3508 1897
<< metal2 >>
rect 3296 1843 3508 1897
<< metal3 >>
rect 3296 1843 3508 1897
<< metal4 >>
rect 3296 1843 3508 1897
<< via3 >>
rect 3303 1850 3501 1890
<< via2 >>
rect 3303 1850 3501 1890
<< via1 >>
rect 3303 1850 3501 1890
<< labels >>
flabel metal3 s 4543 1631 4686 1661 0 FreeSans 400 0 0 0 IN+
port 4 nsew signal bidirectional
flabel metal3 s 3791 831 3934 861 0 FreeSans 400 0 0 0 IN-
port 5 nsew signal bidirectional
flabel metal1 s 0 4056 5600 4106 0 FreeSans 400 0 0 0 VDD
port 6 nsew signal bidirectional
flabel metal1 s 100 3956 5500 4006 0 FreeSans 400 0 0 0 VSS
port 7 nsew signal bidirectional
flabel metal3 s 5073 3296 5232 3326 0 FreeSans 400 0 0 0 OUT
port 8 nsew signal bidirectional
<< properties >>
<< end >>