magic
tech sky130A
magscale 1 1
timestamp 1745832349
<< checkpaint >>
rect 0 0 1 1
use JNWATR_NCH_4C5F0 diff1_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 2260
box 0 0 576 240
use JNWATR_NCH_4C5F0 diff1_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2500
box 0 0 576 400
use JNWATR_NCH_4CTAPBOT diff1_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2260
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 500
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP5_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 260
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 500
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT load1_MP6_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 260
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 1300
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 1700
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 1300
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP load1_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 1700
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror2_MN4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 2900
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror2_MN3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 2900
box 0 0 576 400
use JNWATR_NCH_4C5F0 mirror1_MN5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 3300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN5_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 3700
box 0 0 576 240
use JNWATR_NCH_4C5F0 mirror1_MN6 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 3300
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP mirror1_MN6_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 3700
box 0 0 576 240
use JNWATR_PCH_4C5F0 load1_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 876 0 1 900
box 0 0 576 400
use JNWATR_PCH_4C5F0 load1_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 300 0 1 900
box 0 0 576 400
<< m1 >>
rect 629 513 739 567
<< m2 >>
rect 629 513 739 567
<< m3 >>
rect 629 513 739 567
<< via2 >>
rect 636 520 732 560
<< via1 >>
rect 636 520 732 560
<< m1 >>
rect 629 3313 739 3367
<< m2 >>
rect 629 3313 739 3367
<< m3 >>
rect 629 3313 739 3367
<< via2 >>
rect 636 3320 732 3360
<< via1 >>
rect 636 3320 732 3360
<< m1 >>
rect 373 3073 419 3127
<< m2 >>
rect 373 3073 419 3127
<< via1 >>
rect 380 3080 412 3120
<< m1 >>
rect 373 3073 419 3127
<< m2 >>
rect 373 3073 419 3127
<< m3 >>
rect 373 3073 419 3127
<< via2 >>
rect 380 3080 412 3120
<< via1 >>
rect 380 3080 412 3120
<< m1 >>
rect 949 3073 995 3127
<< m2 >>
rect 949 3073 995 3127
<< m3 >>
rect 949 3073 995 3127
<< via2 >>
rect 956 3080 988 3120
<< via1 >>
rect 956 3080 988 3120
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< m3 >>
rect 1205 2513 1315 2567
<< via2 >>
rect 1212 2520 1308 2560
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< m3 >>
rect 1205 2513 1315 2567
<< via2 >>
rect 1212 2520 1308 2560
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< m3 >>
rect 1205 2513 1315 2567
<< via2 >>
rect 1212 2520 1308 2560
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< m3 >>
rect 373 1473 419 1527
<< via2 >>
rect 380 1480 412 1520
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< m3 >>
rect 373 1473 419 1527
<< via2 >>
rect 380 1480 412 1520
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< m3 >>
rect 949 1473 995 1527
<< via2 >>
rect 956 1480 988 1520
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< m3 >>
rect 949 1473 995 1527
<< via2 >>
rect 956 1480 988 1520
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< m3 >>
rect 1205 1313 1315 1367
<< via2 >>
rect 1212 1320 1308 1360
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< m3 >>
rect 1205 1313 1315 1367
<< via2 >>
rect 1212 1320 1308 1360
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< m3 >>
rect 1205 913 1315 967
<< via2 >>
rect 1212 920 1308 960
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< m3 >>
rect 1205 913 1315 967
<< via2 >>
rect 1212 920 1308 960
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< m3 >>
rect 1205 913 1315 967
<< via2 >>
rect 1212 920 1308 960
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 373 1073 419 1127
<< m2 >>
rect 373 1073 419 1127
<< via1 >>
rect 380 1080 412 1120
<< m1 >>
rect 437 2793 547 2847
<< m2 >>
rect 437 2793 547 2847
<< m3 >>
rect 437 2793 547 2847
<< via2 >>
rect 444 2800 540 2840
<< via1 >>
rect 444 2800 540 2840
<< m1 >>
rect 437 2793 547 2847
<< m2 >>
rect 437 2793 547 2847
<< via1 >>
rect 444 2800 540 2840
<< m1 >>
rect 629 2913 739 2967
<< m2 >>
rect 629 2913 739 2967
<< via1 >>
rect 636 2920 732 2960
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< m3 >>
rect 949 673 995 727
<< via2 >>
rect 956 680 988 720
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< m3 >>
rect 949 673 995 727
<< via2 >>
rect 956 680 988 720
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 373 673 419 727
<< m2 >>
rect 373 673 419 727
<< m3 >>
rect 373 673 419 727
<< via2 >>
rect 380 680 412 720
<< via1 >>
rect 380 680 412 720
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< m3 >>
rect 949 1073 995 1127
<< via2 >>
rect 956 1080 988 1120
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< m3 >>
rect 949 1073 995 1127
<< via2 >>
rect 956 1080 988 1120
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 629 913 739 967
<< m2 >>
rect 629 913 739 967
<< via1 >>
rect 636 920 732 960
<< m1 >>
rect 629 1313 739 1367
<< m2 >>
rect 629 1313 739 1367
<< m3 >>
rect 629 1313 739 1367
<< via2 >>
rect 636 1320 732 1360
<< via1 >>
rect 636 1320 732 1360
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< m3 >>
rect 949 3473 995 3527
<< via2 >>
rect 956 3480 988 3520
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< m3 >>
rect 949 3473 995 3527
<< via2 >>
rect 956 3480 988 3520
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 373 3473 419 3527
<< m2 >>
rect 373 3473 419 3527
<< via1 >>
rect 380 3480 412 3520
<< m3 >>
rect 663 534 693 789
<< m2 >>
rect 663 759 837 789
<< m3 >>
rect 807 759 837 3173
<< m2 >>
rect 663 3143 837 3173
<< m3 >>
rect 663 3143 693 3334
<< m1 >>
rect 629 513 739 567
<< m2 >>
rect 629 513 739 567
<< via1 >>
rect 636 520 732 560
<< m1 >>
rect 629 3313 739 3367
<< m2 >>
rect 629 3313 739 3367
<< via1 >>
rect 636 3320 732 3360
<< m2 >>
rect 656 752 700 796
<< m3 >>
rect 656 752 700 796
<< via2 >>
rect 663 759 693 789
<< m2 >>
rect 800 752 844 796
<< m3 >>
rect 800 752 844 796
<< via2 >>
rect 807 759 837 789
<< m2 >>
rect 800 3136 844 3180
<< m3 >>
rect 800 3136 844 3180
<< via2 >>
rect 807 3143 837 3173
<< m2 >>
rect 656 3136 700 3180
<< m3 >>
rect 656 3136 700 3180
<< via2 >>
rect 663 3143 693 3173
<< m2 >>
rect 215 3079 390 3109
<< m3 >>
rect 215 3079 245 3253
<< m2 >>
rect 215 3223 389 3253
<< m3 >>
rect 359 3047 389 3253
<< m2 >>
rect 359 3047 1413 3077
<< m3 >>
rect 1383 2903 1413 3077
<< m2 >>
rect 1383 2903 1557 2933
<< m3 >>
rect 1527 2903 1557 3157
<< m2 >>
rect 1095 3127 1557 3157
<< m3 >>
rect 1095 2935 1125 3157
<< m2 >>
rect 951 2935 1125 2965
<< m3 >>
rect 951 2935 981 3094
<< m1 >>
rect 373 3073 419 3127
<< m2 >>
rect 373 3073 419 3127
<< via1 >>
rect 380 3080 412 3120
<< m1 >>
rect 373 3073 419 3127
<< m2 >>
rect 373 3073 419 3127
<< via1 >>
rect 380 3080 412 3120
<< m1 >>
rect 949 3073 995 3127
<< m2 >>
rect 949 3073 995 3127
<< via1 >>
rect 956 3080 988 3120
<< m2 >>
rect 208 3072 252 3116
<< m3 >>
rect 208 3072 252 3116
<< via2 >>
rect 215 3079 245 3109
<< m2 >>
rect 208 3216 252 3260
<< m3 >>
rect 208 3216 252 3260
<< via2 >>
rect 215 3223 245 3253
<< m2 >>
rect 352 3216 396 3260
<< m3 >>
rect 352 3216 396 3260
<< via2 >>
rect 359 3223 389 3253
<< m2 >>
rect 352 3040 396 3084
<< m3 >>
rect 352 3040 396 3084
<< via2 >>
rect 359 3047 389 3077
<< m2 >>
rect 1376 3040 1420 3084
<< m3 >>
rect 1376 3040 1420 3084
<< via2 >>
rect 1383 3047 1413 3077
<< m2 >>
rect 1376 2896 1420 2940
<< m3 >>
rect 1376 2896 1420 2940
<< via2 >>
rect 1383 2903 1413 2933
<< m2 >>
rect 1520 2896 1564 2940
<< m3 >>
rect 1520 2896 1564 2940
<< via2 >>
rect 1527 2903 1557 2933
<< m2 >>
rect 1520 3120 1564 3164
<< m3 >>
rect 1520 3120 1564 3164
<< via2 >>
rect 1527 3127 1557 3157
<< m2 >>
rect 1088 3120 1132 3164
<< m3 >>
rect 1088 3120 1132 3164
<< via2 >>
rect 1095 3127 1125 3157
<< m2 >>
rect 1088 2928 1132 2972
<< m3 >>
rect 1088 2928 1132 2972
<< via2 >>
rect 1095 2935 1125 2965
<< m2 >>
rect 944 2928 988 2972
<< m3 >>
rect 944 2928 988 2972
<< via2 >>
rect 951 2935 981 2965
<< m2 >>
rect 235 1083 394 1113
<< m3 >>
rect 235 1083 265 1321
<< m2 >>
rect 235 1291 409 1321
<< m3 >>
rect 379 1291 409 1513
<< m3 >>
rect 379 1483 409 1513
<< m2 >>
rect 379 1483 985 1513
<< m3 >>
rect 955 1483 985 1513
<< m3 >>
rect 955 1291 985 1513
<< m2 >>
rect 955 1291 1273 1321
<< m3 >>
rect 1243 923 1273 1321
<< m3 >>
rect 1243 923 1273 953
<< m2 >>
rect 1243 923 1417 953
<< m3 >>
rect 1387 923 1417 1465
<< m2 >>
rect 1243 1435 1417 1465
<< m3 >>
rect 1243 1435 1273 2553
<< m3 >>
rect 1243 923 1273 2553
<< m2 >>
rect 1243 923 1417 953
<< m3 >>
rect 1387 923 1417 1465
<< m2 >>
rect 1243 1435 1417 1465
<< m3 >>
rect 1243 1435 1273 2538
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 1205 2513 1315 2567
<< m2 >>
rect 1205 2513 1315 2567
<< via1 >>
rect 1212 2520 1308 2560
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 373 1473 419 1527
<< m2 >>
rect 373 1473 419 1527
<< via1 >>
rect 380 1480 412 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 949 1473 995 1527
<< m2 >>
rect 949 1473 995 1527
<< via1 >>
rect 956 1480 988 1520
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 1313 1315 1367
<< m2 >>
rect 1205 1313 1315 1367
<< via1 >>
rect 1212 1320 1308 1360
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 1205 913 1315 967
<< m2 >>
rect 1205 913 1315 967
<< via1 >>
rect 1212 920 1308 960
<< m1 >>
rect 373 1073 419 1127
<< m2 >>
rect 373 1073 419 1127
<< via1 >>
rect 380 1080 412 1120
<< m2 >>
rect 228 1076 272 1120
<< m3 >>
rect 228 1076 272 1120
<< via2 >>
rect 235 1083 265 1113
<< m2 >>
rect 228 1284 272 1328
<< m3 >>
rect 228 1284 272 1328
<< via2 >>
rect 235 1291 265 1321
<< m2 >>
rect 372 1284 416 1328
<< m3 >>
rect 372 1284 416 1328
<< via2 >>
rect 379 1291 409 1321
<< m2 >>
rect 372 1476 416 1520
<< m3 >>
rect 372 1476 416 1520
<< via2 >>
rect 379 1483 409 1513
<< m2 >>
rect 948 1476 992 1520
<< m3 >>
rect 948 1476 992 1520
<< via2 >>
rect 955 1483 985 1513
<< m2 >>
rect 948 1284 992 1328
<< m3 >>
rect 948 1284 992 1328
<< via2 >>
rect 955 1291 985 1321
<< m2 >>
rect 1236 1284 1280 1328
<< m3 >>
rect 1236 1284 1280 1328
<< via2 >>
rect 1243 1291 1273 1321
<< m2 >>
rect 1236 916 1280 960
<< m3 >>
rect 1236 916 1280 960
<< via2 >>
rect 1243 923 1273 953
<< m2 >>
rect 1380 916 1424 960
<< m3 >>
rect 1380 916 1424 960
<< via2 >>
rect 1387 923 1417 953
<< m2 >>
rect 1380 1428 1424 1472
<< m3 >>
rect 1380 1428 1424 1472
<< via2 >>
rect 1387 1435 1417 1465
<< m2 >>
rect 1236 1428 1280 1472
<< m3 >>
rect 1236 1428 1280 1472
<< via2 >>
rect 1243 1435 1273 1465
<< m2 >>
rect 1236 916 1280 960
<< m3 >>
rect 1236 916 1280 960
<< via2 >>
rect 1243 923 1273 953
<< m2 >>
rect 1380 916 1424 960
<< m3 >>
rect 1380 916 1424 960
<< via2 >>
rect 1387 923 1417 953
<< m2 >>
rect 1380 1428 1424 1472
<< m3 >>
rect 1380 1428 1424 1472
<< via2 >>
rect 1387 1435 1417 1465
<< m2 >>
rect 1236 1428 1280 1472
<< m3 >>
rect 1236 1428 1280 1472
<< via2 >>
rect 1243 1435 1273 1465
<< m2 >>
rect 505 2915 680 2945
<< m3 >>
rect 505 2659 535 2945
<< m2 >>
rect 505 2659 679 2689
<< m3 >>
rect 649 2659 679 2833
<< m2 >>
rect 488 2803 679 2833
<< m1 >>
rect 437 2793 547 2847
<< m2 >>
rect 437 2793 547 2847
<< via1 >>
rect 444 2800 540 2840
<< m1 >>
rect 437 2793 547 2847
<< m2 >>
rect 437 2793 547 2847
<< via1 >>
rect 444 2800 540 2840
<< m1 >>
rect 629 2913 739 2967
<< m2 >>
rect 629 2913 739 2967
<< via1 >>
rect 636 2920 732 2960
<< m2 >>
rect 498 2908 542 2952
<< m3 >>
rect 498 2908 542 2952
<< via2 >>
rect 505 2915 535 2945
<< m2 >>
rect 498 2652 542 2696
<< m3 >>
rect 498 2652 542 2696
<< via2 >>
rect 505 2659 535 2689
<< m2 >>
rect 642 2652 686 2696
<< m3 >>
rect 642 2652 686 2696
<< via2 >>
rect 649 2659 679 2689
<< m2 >>
rect 642 2796 686 2840
<< m3 >>
rect 642 2796 686 2840
<< via2 >>
rect 649 2803 679 2833
<< m3 >>
rect 378 411 408 697
<< m2 >>
rect 378 411 984 441
<< m3 >>
rect 954 411 984 712
<< m3 >>
rect 954 682 984 712
<< m2 >>
rect 954 682 1512 712
<< m3 >>
rect 1482 682 1512 1112
<< m2 >>
rect 954 1082 1512 1112
<< m3 >>
rect 954 1082 984 1112
<< m3 >>
rect 954 922 984 1112
<< m2 >>
rect 681 922 984 952
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 949 673 995 727
<< m2 >>
rect 949 673 995 727
<< via1 >>
rect 956 680 988 720
<< m1 >>
rect 373 673 419 727
<< m2 >>
rect 373 673 419 727
<< via1 >>
rect 380 680 412 720
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 949 1073 995 1127
<< m2 >>
rect 949 1073 995 1127
<< via1 >>
rect 956 1080 988 1120
<< m1 >>
rect 629 913 739 967
<< m2 >>
rect 629 913 739 967
<< via1 >>
rect 636 920 732 960
<< m2 >>
rect 371 404 415 448
<< m3 >>
rect 371 404 415 448
<< via2 >>
rect 378 411 408 441
<< m2 >>
rect 947 404 991 448
<< m3 >>
rect 947 404 991 448
<< via2 >>
rect 954 411 984 441
<< m2 >>
rect 947 675 991 719
<< m3 >>
rect 947 675 991 719
<< via2 >>
rect 954 682 984 712
<< m2 >>
rect 1475 675 1519 719
<< m3 >>
rect 1475 675 1519 719
<< via2 >>
rect 1482 682 1512 712
<< m2 >>
rect 1475 1075 1519 1119
<< m3 >>
rect 1475 1075 1519 1119
<< via2 >>
rect 1482 1082 1512 1112
<< m2 >>
rect 947 1075 991 1119
<< m3 >>
rect 947 1075 991 1119
<< via2 >>
rect 954 1082 984 1112
<< m2 >>
rect 947 915 991 959
<< m3 >>
rect 947 915 991 959
<< via2 >>
rect 954 922 984 952
<< m2 >>
rect 392 3481 983 3511
<< m3 >>
rect 953 3481 983 3511
<< m3 >>
rect 953 3337 983 3511
<< m2 >>
rect 953 3337 1127 3367
<< m3 >>
rect 1097 3337 1127 3511
<< m2 >>
rect 1097 3481 1511 3511
<< m3 >>
rect 1481 3337 1511 3511
<< m2 >>
rect 1481 3337 1655 3367
<< m3 >>
rect 1625 2697 1655 3367
<< m2 >>
rect 1465 2697 1655 2727
<< m3 >>
rect 1465 2169 1495 2727
<< m2 >>
rect 1145 2169 1495 2199
<< m3 >>
rect 1145 1881 1175 2199
<< m2 >>
rect 1001 1881 1175 1911
<< m3 >>
rect 1001 1721 1031 1911
<< m2 >>
rect 665 1721 1031 1751
<< m3 >>
rect 665 1336 695 1751
<< m1 >>
rect 629 1313 739 1367
<< m2 >>
rect 629 1313 739 1367
<< via1 >>
rect 636 1320 732 1360
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 949 3473 995 3527
<< m2 >>
rect 949 3473 995 3527
<< via1 >>
rect 956 3480 988 3520
<< m1 >>
rect 373 3473 419 3527
<< m2 >>
rect 373 3473 419 3527
<< via1 >>
rect 380 3480 412 3520
<< m2 >>
rect 946 3474 990 3518
<< m3 >>
rect 946 3474 990 3518
<< via2 >>
rect 953 3481 983 3511
<< m2 >>
rect 946 3330 990 3374
<< m3 >>
rect 946 3330 990 3374
<< via2 >>
rect 953 3337 983 3367
<< m2 >>
rect 1090 3330 1134 3374
<< m3 >>
rect 1090 3330 1134 3374
<< via2 >>
rect 1097 3337 1127 3367
<< m2 >>
rect 1090 3474 1134 3518
<< m3 >>
rect 1090 3474 1134 3518
<< via2 >>
rect 1097 3481 1127 3511
<< m2 >>
rect 1474 3474 1518 3518
<< m3 >>
rect 1474 3474 1518 3518
<< via2 >>
rect 1481 3481 1511 3511
<< m2 >>
rect 1474 3330 1518 3374
<< m3 >>
rect 1474 3330 1518 3374
<< via2 >>
rect 1481 3337 1511 3367
<< m2 >>
rect 1618 3330 1662 3374
<< m3 >>
rect 1618 3330 1662 3374
<< via2 >>
rect 1625 3337 1655 3367
<< m2 >>
rect 1618 2690 1662 2734
<< m3 >>
rect 1618 2690 1662 2734
<< via2 >>
rect 1625 2697 1655 2727
<< m2 >>
rect 1458 2690 1502 2734
<< m3 >>
rect 1458 2690 1502 2734
<< via2 >>
rect 1465 2697 1495 2727
<< m2 >>
rect 1458 2162 1502 2206
<< m3 >>
rect 1458 2162 1502 2206
<< via2 >>
rect 1465 2169 1495 2199
<< m2 >>
rect 1138 2162 1182 2206
<< m3 >>
rect 1138 2162 1182 2206
<< via2 >>
rect 1145 2169 1175 2199
<< m2 >>
rect 1138 1874 1182 1918
<< m3 >>
rect 1138 1874 1182 1918
<< via2 >>
rect 1145 1881 1175 1911
<< m2 >>
rect 994 1874 1038 1918
<< m3 >>
rect 994 1874 1038 1918
<< via2 >>
rect 1001 1881 1031 1911
<< m2 >>
rect 994 1714 1038 1758
<< m3 >>
rect 994 1714 1038 1758
<< via2 >>
rect 1001 1721 1031 1751
<< m2 >>
rect 658 1714 702 1758
<< m3 >>
rect 658 1714 702 1758
<< via2 >>
rect 665 1721 695 1751
<< locali >>
rect 100 4050 1652 4100
<< locali >>
rect 100 100 1652 150
<< m1 >>
rect 100 150 150 4050
<< m1 >>
rect 1602 150 1652 4050
<< locali >>
rect 93 4043 157 4107
<< m1 >>
rect 93 4043 157 4107
<< viali >>
rect 100 4050 150 4100
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1595 4043 1659 4107
<< m1 >>
rect 1595 4043 1659 4107
<< viali >>
rect 1602 4050 1652 4100
<< locali >>
rect 1595 93 1659 157
<< m1 >>
rect 1595 93 1659 157
<< viali >>
rect 1602 100 1652 150
<< locali >>
rect 0 4150 1752 4200
<< locali >>
rect 0 0 1752 50
<< m1 >>
rect 0 50 50 4150
<< m1 >>
rect 1702 50 1752 4150
<< locali >>
rect -7 4143 57 4207
<< m1 >>
rect -7 4143 57 4207
<< viali >>
rect 0 4150 50 4200
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1695 4143 1759 4207
<< m1 >>
rect 1695 4143 1759 4207
<< viali >>
rect 1702 4150 1752 4200
<< locali >>
rect 1695 -7 1759 57
<< m1 >>
rect 1695 -7 1759 57
<< viali >>
rect 1702 0 1752 50
<< locali >>
rect 828 800 1116 840
<< locali >>
rect 1212 680 1372 720
<< locali >>
rect 252 800 540 840
<< locali >>
rect 252 1600 540 1640
<< locali >>
rect 828 1600 1116 1640
<< locali >>
rect 1212 1480 1372 1520
<< locali >>
rect 252 3200 540 3240
<< locali >>
rect 828 3200 1116 3240
<< locali >>
rect 1212 3080 1372 3120
<< locali >>
rect 828 3600 1116 3640
<< locali >>
rect 1212 3480 1372 3520
<< locali >>
rect 252 3600 540 3640
<< locali >>
rect 828 1200 1116 1240
<< locali >>
rect 252 1200 540 1240
<< locali >>
rect 0 2332 1752 2428
<< locali >>
rect -7 2325 57 2435
<< m1 >>
rect -7 2325 57 2435
<< viali >>
rect 0 2332 50 2428
<< locali >>
rect 1695 2325 1759 2435
<< m1 >>
rect 1695 2325 1759 2435
<< viali >>
rect 1702 2332 1752 2428
<< locali >>
rect 100 332 1652 428
<< locali >>
rect 93 325 157 435
<< m1 >>
rect 93 325 157 435
<< viali >>
rect 100 332 150 428
<< locali >>
rect 1595 325 1659 435
<< m1 >>
rect 1595 325 1659 435
<< viali >>
rect 1602 332 1652 428
<< locali >>
rect 100 1772 1652 1868
<< locali >>
rect 93 1765 157 1875
<< m1 >>
rect 93 1765 157 1875
<< viali >>
rect 100 1772 150 1868
<< locali >>
rect 1595 1765 1659 1875
<< m1 >>
rect 1595 1765 1659 1875
<< viali >>
rect 1602 1772 1652 1868
<< locali >>
rect 0 3772 1752 3868
<< locali >>
rect -7 3765 57 3875
<< m1 >>
rect -7 3765 57 3875
<< viali >>
rect 0 3772 50 3868
<< locali >>
rect 1695 3765 1759 3875
<< m1 >>
rect 1695 3765 1759 3875
<< viali >>
rect 1702 3772 1752 3868
<< labels >>
flabel locali s 0 4150 1752 4200 0 FreeSans 400 0 0 0 VSS
port 327 nsew signal bidirectional
flabel locali s 100 4050 1652 4100 0 FreeSans 400 0 0 0 VDD
port 328 nsew signal bidirectional
flabel m1 s 956 2680 988 2720 0 FreeSans 400 0 0 0 VIP
port 329 nsew signal bidirectional
flabel m1 s 380 2680 412 2720 0 FreeSans 400 0 0 0 VIN
port 330 nsew signal bidirectional
flabel m3 s 663 534 693 789 0 FreeSans 400 0 0 0 VO
port 331 nsew signal bidirectional
flabel m2 s 215 3079 390 3109 0 FreeSans 400 0 0 0 I_BIAS
port 332 nsew signal bidirectional
<< properties >>
<< end >>