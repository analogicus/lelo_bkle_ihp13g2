magic
tech sky130A
magscale 1 1
timestamp 1746459945
<< checkpaint >>
rect 0 0 1 1
use JNWATR_PCH_4C5F0 None_MP2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 2600
box 0 0 576 240
use JNWATR_PCH_4CTAPBOT None_MP2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1960
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2200
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 2600
box 0 0 576 240
use AALMISC_CAP50f None_CM1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 2646
box 0 0 580 842
use JNWATR_PCH_4C5F0 None_MP3 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPTOP None_MP3_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1800
box 0 0 576 240
use JNWATR_PCH_4CTAPBOT None_MP3_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP4 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1400
box 0 0 576 400
use JNWATR_PCH_4CTAPBOT None_MP4_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1160
box 0 0 576 240
use JNWATR_PCH_4C5F0 None_MP5 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 1800
box 0 0 576 400
use JNWATR_NCH_4C5F0 None_MN1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN1_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN1_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 292 0 1 -40
box 0 0 576 240
use JNWATR_NCH_4C5F0 None_MN2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 200
box 0 0 576 400
use JNWATR_NCH_4CTAPTOP None_MN2_TAPTOP ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 600
box 0 0 576 240
use JNWATR_NCH_4CTAPBOT None_MN2_TAPBOT ~/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A
transform 1 0 868 0 1 -40
box 0 0 576 240
use JNWTR_RPPO8 None_RH2 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 3838
box 0 0 1372 1720
use JNWTR_RPPO4 None_RH1 ~/aicex/ip/jnw_bkle_sky130A/design/JNW_TR_SKY130A
transform 1 0 200 0 1 5608
box 0 0 940 1720
use AALMISC_PNP_W3p40L3p40 load1_QP1 ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 13438
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<0> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 9118
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<1> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 10558
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<2> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 9838
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<3> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 12718
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<4> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 7678
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<5> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 11998
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<6> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 8398
box 0 0 670 670
use AALMISC_PNP_W3p40L3p40 load1_QP2<7> ~/aicex/ip/jnw_bkle_sky130A/design/AAL_MISC_SKY130A
transform 1 0 200 0 1 11278
box 0 0 670 670
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< m3 >>
rect 621 2213 731 2267
<< via2 >>
rect 628 2220 724 2260
<< via1 >>
rect 628 2220 724 2260
<< locali >>
rect 375 7061 533 7195
<< m1 >>
rect 375 7061 533 7195
<< m2 >>
rect 375 7061 533 7195
<< m3 >>
rect 375 7061 533 7195
<< via2 >>
rect 382 7068 526 7188
<< via1 >>
rect 382 7068 526 7188
<< viali >>
rect 382 7068 526 7188
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< m3 >>
rect 365 2373 411 2427
<< via2 >>
rect 372 2380 404 2420
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< m3 >>
rect 941 2373 987 2427
<< via2 >>
rect 948 2380 980 2420
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m1 >>
rect 1197 2213 1307 2267
<< m2 >>
rect 1197 2213 1307 2267
<< m3 >>
rect 1197 2213 1307 2267
<< via2 >>
rect 1204 2220 1300 2260
<< via1 >>
rect 1204 2220 1300 2260
<< m1 >>
rect 463 13744 607 13810
<< m2 >>
rect 463 13744 607 13810
<< via1 >>
rect 470 13751 600 13803
<< m1 >>
rect 621 1413 731 1467
<< m2 >>
rect 621 1413 731 1467
<< m3 >>
rect 621 1413 731 1467
<< via2 >>
rect 628 1420 724 1460
<< via1 >>
rect 628 1420 724 1460
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< m3 >>
rect 621 213 731 267
<< via2 >>
rect 628 220 724 260
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< m3 >>
rect 621 213 731 267
<< via2 >>
rect 628 220 724 260
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< m3 >>
rect 621 213 731 267
<< via2 >>
rect 628 220 724 260
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< m3 >>
rect 941 1573 987 1627
<< via2 >>
rect 948 1580 980 1620
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< m3 >>
rect 1197 1413 1307 1467
<< via2 >>
rect 1204 1420 1300 1460
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 941 1973 987 2027
<< m2 >>
rect 941 1973 987 2027
<< via1 >>
rect 948 1980 980 2020
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< m3 >>
rect 1197 213 1307 267
<< via2 >>
rect 1204 220 1300 260
<< via1 >>
rect 1204 220 1300 260
<< locali >>
rect 375 5291 533 5425
<< m1 >>
rect 375 5291 533 5425
<< m2 >>
rect 375 5291 533 5425
<< via1 >>
rect 382 5298 526 5418
<< viali >>
rect 382 5298 526 5418
<< locali >>
rect 807 7061 965 7195
<< m1 >>
rect 807 7061 965 7195
<< m2 >>
rect 807 7061 965 7195
<< via1 >>
rect 814 7068 958 7188
<< viali >>
rect 814 7068 958 7188
<< locali >>
rect 1239 5291 1397 5425
<< m1 >>
rect 1239 5291 1397 5425
<< m2 >>
rect 1239 5291 1397 5425
<< m3 >>
rect 1239 5291 1397 5425
<< via2 >>
rect 1246 5298 1390 5418
<< via1 >>
rect 1246 5298 1390 5418
<< viali >>
rect 1246 5298 1390 5418
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< m3 >>
rect 463 9424 607 9490
<< via2 >>
rect 470 9431 600 9483
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< m3 >>
rect 463 10864 607 10930
<< via2 >>
rect 470 10871 600 10923
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< m3 >>
rect 463 10144 607 10210
<< via2 >>
rect 470 10151 600 10203
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 13024 607 13090
<< m2 >>
rect 463 13024 607 13090
<< via1 >>
rect 470 13031 600 13083
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< m3 >>
rect 463 7984 607 8050
<< via2 >>
rect 470 7991 600 8043
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< m3 >>
rect 463 12304 607 12370
<< via2 >>
rect 470 12311 600 12363
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< m3 >>
rect 463 8704 607 8770
<< via2 >>
rect 470 8711 600 8763
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< via1 >>
rect 470 11591 600 11643
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< m3 >>
rect 463 11584 607 11650
<< via2 >>
rect 470 11591 600 11643
<< via1 >>
rect 470 11591 600 11643
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< via1 >>
rect 470 11591 600 11643
<< m3 >>
rect 657 2234 687 2697
<< m2 >>
rect 657 2667 879 2697
<< m3 >>
rect 849 2667 879 6985
<< m2 >>
rect 433 6955 879 6985
<< m3 >>
rect 433 6955 463 7130
<< m1 >>
rect 621 2213 731 2267
<< m2 >>
rect 621 2213 731 2267
<< via1 >>
rect 628 2220 724 2260
<< locali >>
rect 375 7061 533 7195
<< m1 >>
rect 375 7061 533 7195
<< viali >>
rect 382 7068 526 7188
<< m2 >>
rect 650 2660 694 2704
<< m3 >>
rect 650 2660 694 2704
<< via2 >>
rect 657 2667 687 2697
<< m2 >>
rect 842 2660 886 2704
<< m3 >>
rect 842 2660 886 2704
<< via2 >>
rect 849 2667 879 2697
<< m2 >>
rect 842 6948 886 6992
<< m3 >>
rect 842 6948 886 6992
<< via2 >>
rect 849 6955 879 6985
<< m2 >>
rect 426 6948 470 6992
<< m3 >>
rect 426 6948 470 6992
<< via2 >>
rect 433 6955 463 6985
<< m2 >>
rect 245 1583 388 1613
<< m3 >>
rect 245 1583 275 2413
<< m2 >>
rect 245 2383 403 2413
<< m3 >>
rect 373 2383 403 2413
<< m2 >>
rect 373 2383 979 2413
<< m3 >>
rect 949 2383 979 2413
<< m2 >>
rect 341 2383 979 2413
<< m3 >>
rect 341 2383 371 2717
<< m2 >>
rect 341 2687 484 2717
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 365 2373 411 2427
<< m2 >>
rect 365 2373 411 2427
<< via1 >>
rect 372 2380 404 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 941 2373 987 2427
<< m2 >>
rect 941 2373 987 2427
<< via1 >>
rect 948 2380 980 2420
<< m1 >>
rect 365 1573 411 1627
<< m2 >>
rect 365 1573 411 1627
<< via1 >>
rect 372 1580 404 1620
<< m2 >>
rect 238 1576 282 1620
<< m3 >>
rect 238 1576 282 1620
<< via2 >>
rect 245 1583 275 1613
<< m2 >>
rect 238 2376 282 2420
<< m3 >>
rect 238 2376 282 2420
<< via2 >>
rect 245 2383 275 2413
<< m2 >>
rect 366 2376 410 2420
<< m3 >>
rect 366 2376 410 2420
<< via2 >>
rect 373 2383 403 2413
<< m2 >>
rect 366 2376 410 2420
<< m3 >>
rect 366 2376 410 2420
<< via2 >>
rect 373 2383 403 2413
<< m2 >>
rect 942 2376 986 2420
<< m3 >>
rect 942 2376 986 2420
<< via2 >>
rect 949 2383 979 2413
<< m2 >>
rect 942 2376 986 2420
<< m3 >>
rect 942 2376 986 2420
<< via2 >>
rect 949 2383 979 2413
<< m2 >>
rect 334 2376 378 2420
<< m3 >>
rect 334 2376 378 2420
<< via2 >>
rect 341 2383 371 2413
<< m2 >>
rect 334 2680 378 2724
<< m3 >>
rect 334 2680 378 2724
<< via2 >>
rect 341 2687 371 2717
<< m3 >>
rect 1233 2234 1263 5209
<< m2 >>
rect 689 5179 1263 5209
<< m3 >>
rect 689 5179 719 13785
<< m2 >>
rect 528 13755 719 13785
<< m1 >>
rect 1197 2213 1307 2267
<< m2 >>
rect 1197 2213 1307 2267
<< via1 >>
rect 1204 2220 1300 2260
<< m1 >>
rect 463 13744 607 13810
<< m2 >>
rect 463 13744 607 13810
<< via1 >>
rect 470 13751 600 13803
<< m2 >>
rect 1226 5172 1270 5216
<< m3 >>
rect 1226 5172 1270 5216
<< via2 >>
rect 1233 5179 1263 5209
<< m2 >>
rect 682 5172 726 5216
<< m3 >>
rect 682 5172 726 5216
<< via2 >>
rect 689 5179 719 5209
<< m2 >>
rect 682 13748 726 13792
<< m3 >>
rect 682 13748 726 13792
<< via2 >>
rect 689 13755 719 13785
<< m2 >>
rect 658 381 961 411
<< m3 >>
rect 658 221 688 411
<< m3 >>
rect 658 221 688 251
<< m3 >>
rect 658 221 688 1436
<< m1 >>
rect 621 1413 731 1467
<< m2 >>
rect 621 1413 731 1467
<< via1 >>
rect 628 1420 724 1460
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 621 213 731 267
<< m2 >>
rect 621 213 731 267
<< via1 >>
rect 628 220 724 260
<< m1 >>
rect 941 373 987 427
<< m2 >>
rect 941 373 987 427
<< via1 >>
rect 948 380 980 420
<< m2 >>
rect 651 374 695 418
<< m3 >>
rect 651 374 695 418
<< via2 >>
rect 658 381 688 411
<< m3 >>
rect 1235 237 1265 1452
<< m3 >>
rect 1235 1422 1265 1452
<< m3 >>
rect 1235 1422 1265 1612
<< m2 >>
rect 947 1582 1265 1612
<< m3 >>
rect 947 1582 977 1612
<< m2 >>
rect 819 1582 977 1612
<< m3 >>
rect 819 1582 849 2012
<< m2 >>
rect 819 1982 962 2012
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 941 1573 987 1627
<< m2 >>
rect 941 1573 987 1627
<< via1 >>
rect 948 1580 980 1620
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 1197 1413 1307 1467
<< m2 >>
rect 1197 1413 1307 1467
<< via1 >>
rect 1204 1420 1300 1460
<< m1 >>
rect 941 1973 987 2027
<< m2 >>
rect 941 1973 987 2027
<< via1 >>
rect 948 1980 980 2020
<< m1 >>
rect 1197 213 1307 267
<< m2 >>
rect 1197 213 1307 267
<< via1 >>
rect 1204 220 1300 260
<< m2 >>
rect 1228 1575 1272 1619
<< m3 >>
rect 1228 1575 1272 1619
<< via2 >>
rect 1235 1582 1265 1612
<< m2 >>
rect 940 1575 984 1619
<< m3 >>
rect 940 1575 984 1619
<< via2 >>
rect 947 1582 977 1612
<< m2 >>
rect 940 1575 984 1619
<< m3 >>
rect 940 1575 984 1619
<< via2 >>
rect 947 1582 977 1612
<< m2 >>
rect 812 1575 856 1619
<< m3 >>
rect 812 1575 856 1619
<< via2 >>
rect 819 1582 849 1612
<< m2 >>
rect 812 1975 856 2019
<< m3 >>
rect 812 1975 856 2019
<< via2 >>
rect 819 1982 849 2012
<< m2 >>
rect 449 5338 624 5368
<< m3 >>
rect 594 5338 624 7144
<< m2 >>
rect 594 7114 881 7144
<< locali >>
rect 375 5291 533 5425
<< m1 >>
rect 375 5291 533 5425
<< viali >>
rect 382 5298 526 5418
<< locali >>
rect 807 7061 965 7195
<< m1 >>
rect 807 7061 965 7195
<< viali >>
rect 814 7068 958 7188
<< m2 >>
rect 587 5331 631 5375
<< m3 >>
rect 587 5331 631 5375
<< via2 >>
rect 594 5338 624 5368
<< m2 >>
rect 587 7107 631 7151
<< m3 >>
rect 587 7107 631 7151
<< via2 >>
rect 594 7114 624 7144
<< m2 >>
rect 391 13040 534 13070
<< m3 >>
rect 391 12320 421 13070
<< m2 >>
rect 391 12320 549 12350
<< m3 >>
rect 519 12320 549 12350
<< m2 >>
rect 391 12320 549 12350
<< m3 >>
rect 391 11600 421 12350
<< m2 >>
rect 391 11600 549 11630
<< m3 >>
rect 519 11600 549 11630
<< m2 >>
rect 391 11600 549 11630
<< m3 >>
rect 391 10880 421 11630
<< m2 >>
rect 391 10880 549 10910
<< m3 >>
rect 519 10880 549 10910
<< m2 >>
rect 391 10880 549 10910
<< m3 >>
rect 391 10160 421 10910
<< m2 >>
rect 391 10160 549 10190
<< m3 >>
rect 519 10160 549 10190
<< m2 >>
rect 391 10160 549 10190
<< m3 >>
rect 391 9440 421 10190
<< m2 >>
rect 391 9440 549 9470
<< m3 >>
rect 519 9440 549 9470
<< m2 >>
rect 391 9440 549 9470
<< m3 >>
rect 391 8720 421 9470
<< m2 >>
rect 391 8720 549 8750
<< m3 >>
rect 519 8720 549 8750
<< m2 >>
rect 391 8720 549 8750
<< m3 >>
rect 391 8000 421 8750
<< m2 >>
rect 391 8000 549 8030
<< m3 >>
rect 519 8000 549 8030
<< m2 >>
rect 519 8000 1333 8030
<< m3 >>
rect 1303 5359 1333 8030
<< locali >>
rect 1239 5291 1397 5425
<< m1 >>
rect 1239 5291 1397 5425
<< viali >>
rect 1246 5298 1390 5418
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 9424 607 9490
<< m2 >>
rect 463 9424 607 9490
<< via1 >>
rect 470 9431 600 9483
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10864 607 10930
<< m2 >>
rect 463 10864 607 10930
<< via1 >>
rect 470 10871 600 10923
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 10144 607 10210
<< m2 >>
rect 463 10144 607 10210
<< via1 >>
rect 470 10151 600 10203
<< m1 >>
rect 463 13024 607 13090
<< m2 >>
rect 463 13024 607 13090
<< via1 >>
rect 470 13031 600 13083
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 7984 607 8050
<< m2 >>
rect 463 7984 607 8050
<< via1 >>
rect 470 7991 600 8043
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 12304 607 12370
<< m2 >>
rect 463 12304 607 12370
<< via1 >>
rect 470 12311 600 12363
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 8704 607 8770
<< m2 >>
rect 463 8704 607 8770
<< via1 >>
rect 470 8711 600 8763
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< via1 >>
rect 470 11591 600 11643
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< via1 >>
rect 470 11591 600 11643
<< m1 >>
rect 463 11584 607 11650
<< m2 >>
rect 463 11584 607 11650
<< via1 >>
rect 470 11591 600 11643
<< m2 >>
rect 384 13033 428 13077
<< m3 >>
rect 384 13033 428 13077
<< via2 >>
rect 391 13040 421 13070
<< m2 >>
rect 384 12313 428 12357
<< m3 >>
rect 384 12313 428 12357
<< via2 >>
rect 391 12320 421 12350
<< m2 >>
rect 512 12313 556 12357
<< m3 >>
rect 512 12313 556 12357
<< via2 >>
rect 519 12320 549 12350
<< m2 >>
rect 512 12313 556 12357
<< m3 >>
rect 512 12313 556 12357
<< via2 >>
rect 519 12320 549 12350
<< m2 >>
rect 384 12313 428 12357
<< m3 >>
rect 384 12313 428 12357
<< via2 >>
rect 391 12320 421 12350
<< m2 >>
rect 384 11593 428 11637
<< m3 >>
rect 384 11593 428 11637
<< via2 >>
rect 391 11600 421 11630
<< m2 >>
rect 512 11593 556 11637
<< m3 >>
rect 512 11593 556 11637
<< via2 >>
rect 519 11600 549 11630
<< m2 >>
rect 512 11593 556 11637
<< m3 >>
rect 512 11593 556 11637
<< via2 >>
rect 519 11600 549 11630
<< m2 >>
rect 384 11593 428 11637
<< m3 >>
rect 384 11593 428 11637
<< via2 >>
rect 391 11600 421 11630
<< m2 >>
rect 384 10873 428 10917
<< m3 >>
rect 384 10873 428 10917
<< via2 >>
rect 391 10880 421 10910
<< m2 >>
rect 512 10873 556 10917
<< m3 >>
rect 512 10873 556 10917
<< via2 >>
rect 519 10880 549 10910
<< m2 >>
rect 512 10873 556 10917
<< m3 >>
rect 512 10873 556 10917
<< via2 >>
rect 519 10880 549 10910
<< m2 >>
rect 384 10873 428 10917
<< m3 >>
rect 384 10873 428 10917
<< via2 >>
rect 391 10880 421 10910
<< m2 >>
rect 384 10153 428 10197
<< m3 >>
rect 384 10153 428 10197
<< via2 >>
rect 391 10160 421 10190
<< m2 >>
rect 512 10153 556 10197
<< m3 >>
rect 512 10153 556 10197
<< via2 >>
rect 519 10160 549 10190
<< m2 >>
rect 512 10153 556 10197
<< m3 >>
rect 512 10153 556 10197
<< via2 >>
rect 519 10160 549 10190
<< m2 >>
rect 384 10153 428 10197
<< m3 >>
rect 384 10153 428 10197
<< via2 >>
rect 391 10160 421 10190
<< m2 >>
rect 384 9433 428 9477
<< m3 >>
rect 384 9433 428 9477
<< via2 >>
rect 391 9440 421 9470
<< m2 >>
rect 512 9433 556 9477
<< m3 >>
rect 512 9433 556 9477
<< via2 >>
rect 519 9440 549 9470
<< m2 >>
rect 512 9433 556 9477
<< m3 >>
rect 512 9433 556 9477
<< via2 >>
rect 519 9440 549 9470
<< m2 >>
rect 384 9433 428 9477
<< m3 >>
rect 384 9433 428 9477
<< via2 >>
rect 391 9440 421 9470
<< m2 >>
rect 384 8713 428 8757
<< m3 >>
rect 384 8713 428 8757
<< via2 >>
rect 391 8720 421 8750
<< m2 >>
rect 512 8713 556 8757
<< m3 >>
rect 512 8713 556 8757
<< via2 >>
rect 519 8720 549 8750
<< m2 >>
rect 512 8713 556 8757
<< m3 >>
rect 512 8713 556 8757
<< via2 >>
rect 519 8720 549 8750
<< m2 >>
rect 384 8713 428 8757
<< m3 >>
rect 384 8713 428 8757
<< via2 >>
rect 391 8720 421 8750
<< m2 >>
rect 384 7993 428 8037
<< m3 >>
rect 384 7993 428 8037
<< via2 >>
rect 391 8000 421 8030
<< m2 >>
rect 512 7993 556 8037
<< m3 >>
rect 512 7993 556 8037
<< via2 >>
rect 519 8000 549 8030
<< m2 >>
rect 512 7993 556 8037
<< m3 >>
rect 512 7993 556 8037
<< via2 >>
rect 519 8000 549 8030
<< m2 >>
rect 1296 7993 1340 8037
<< m3 >>
rect 1296 7993 1340 8037
<< via2 >>
rect 1303 8000 1333 8030
<< locali >>
rect 100 14158 1672 14208
<< locali >>
rect 100 100 1672 150
<< m1 >>
rect 100 150 150 14158
<< m1 >>
rect 1622 150 1672 14158
<< locali >>
rect 93 14151 157 14215
<< m1 >>
rect 93 14151 157 14215
<< viali >>
rect 100 14158 150 14208
<< locali >>
rect 93 93 157 157
<< m1 >>
rect 93 93 157 157
<< viali >>
rect 100 100 150 150
<< locali >>
rect 1615 14151 1679 14215
<< m1 >>
rect 1615 14151 1679 14215
<< viali >>
rect 1622 14158 1672 14208
<< locali >>
rect 1615 93 1679 157
<< m1 >>
rect 1615 93 1679 157
<< viali >>
rect 1622 100 1672 150
<< locali >>
rect 0 14258 1772 14308
<< locali >>
rect 0 0 1772 50
<< m1 >>
rect 0 50 50 14258
<< m1 >>
rect 1722 50 1772 14258
<< locali >>
rect -7 14251 57 14315
<< m1 >>
rect -7 14251 57 14315
<< viali >>
rect 0 14258 50 14308
<< locali >>
rect -7 -7 57 57
<< m1 >>
rect -7 -7 57 57
<< viali >>
rect 0 0 50 50
<< locali >>
rect 1715 14251 1779 14315
<< m1 >>
rect 1715 14251 1779 14315
<< viali >>
rect 1722 14258 1772 14308
<< locali >>
rect 1715 -7 1779 57
<< m1 >>
rect 1715 -7 1779 57
<< viali >>
rect 1722 0 1772 50
<< locali >>
rect 100 5502 1672 5558
<< locali >>
rect 93 5495 157 5565
<< m1 >>
rect 93 5495 157 5565
<< viali >>
rect 100 5502 150 5558
<< locali >>
rect 1615 5495 1679 5565
<< m1 >>
rect 1615 5495 1679 5565
<< viali >>
rect 1622 5502 1672 5558
<< locali >>
rect 100 3838 1672 3894
<< locali >>
rect 93 3831 157 3901
<< m1 >>
rect 93 3831 157 3901
<< viali >>
rect 100 3838 150 3894
<< locali >>
rect 1615 3831 1679 3901
<< m1 >>
rect 1615 3831 1679 3901
<< viali >>
rect 1622 3838 1672 3894
<< locali >>
rect 100 7272 1672 7328
<< locali >>
rect 93 7265 157 7335
<< m1 >>
rect 93 7265 157 7335
<< viali >>
rect 100 7272 150 7328
<< locali >>
rect 1615 7265 1679 7335
<< m1 >>
rect 1615 7265 1679 7335
<< viali >>
rect 1622 7272 1672 7328
<< locali >>
rect 100 5608 1672 5664
<< locali >>
rect 93 5601 157 5671
<< m1 >>
rect 93 5601 157 5671
<< viali >>
rect 100 5608 150 5664
<< locali >>
rect 1615 5601 1679 5671
<< m1 >>
rect 1615 5601 1679 5671
<< viali >>
rect 1622 5608 1672 5664
<< locali >>
rect 244 2500 532 2540
<< locali >>
rect 820 2500 1108 2540
<< locali >>
rect 244 1700 532 1740
<< locali >>
rect 820 1700 1108 1740
<< locali >>
rect 1204 1580 1364 1620
<< locali >>
rect 820 2100 1108 2140
<< locali >>
rect 244 500 532 540
<< locali >>
rect 628 380 788 420
<< locali >>
rect 820 500 1108 540
<< locali >>
rect 0 2672 1772 2768
<< locali >>
rect -7 2665 57 2775
<< m1 >>
rect -7 2665 57 2775
<< viali >>
rect 0 2672 50 2768
<< locali >>
rect 1715 2665 1779 2775
<< m1 >>
rect 1715 2665 1779 2775
<< viali >>
rect 1722 2672 1772 2768
<< locali >>
rect 0 1232 1772 1328
<< locali >>
rect -7 1225 57 1335
<< m1 >>
rect -7 1225 57 1335
<< viali >>
rect 0 1232 50 1328
<< locali >>
rect 1715 1225 1779 1335
<< m1 >>
rect 1715 1225 1779 1335
<< viali >>
rect 1722 1232 1772 1328
<< locali >>
rect 100 672 1672 768
<< locali >>
rect 93 665 157 775
<< m1 >>
rect 93 665 157 775
<< viali >>
rect 100 672 150 768
<< locali >>
rect 1615 665 1679 775
<< m1 >>
rect 1615 665 1679 775
<< viali >>
rect 1622 672 1672 768
<< locali >>
rect 100 32 1672 128
<< locali >>
rect 93 25 157 135
<< m1 >>
rect 93 25 157 135
<< viali >>
rect 100 32 150 128
<< locali >>
rect 1615 25 1679 135
<< m1 >>
rect 1615 25 1679 135
<< viali >>
rect 1622 32 1672 128
<< locali >>
rect 510 14013 560 14046
<< locali >>
rect 510 9693 560 9726
<< locali >>
rect 510 11133 560 11166
<< locali >>
rect 510 10413 560 10446
<< locali >>
rect 510 13293 560 13326
<< locali >>
rect 510 8253 560 8286
<< locali >>
rect 510 12573 560 12606
<< locali >>
rect 510 8973 560 9006
<< locali >>
rect 510 11853 560 11886
<< locali >>
rect 100 14059 1672 14108
<< locali >>
rect 93 14052 157 14115
<< m1 >>
rect 93 14052 157 14115
<< viali >>
rect 100 14059 150 14108
<< locali >>
rect 1615 14052 1679 14115
<< m1 >>
rect 1615 14052 1679 14115
<< viali >>
rect 1622 14059 1672 14108
<< locali >>
rect 100 13438 1672 13487
<< locali >>
rect 93 13431 157 13494
<< m1 >>
rect 93 13431 157 13494
<< viali >>
rect 100 13438 150 13487
<< locali >>
rect 1615 13431 1679 13494
<< m1 >>
rect 1615 13431 1679 13494
<< viali >>
rect 1622 13438 1672 13487
<< locali >>
rect 100 9739 1672 9788
<< locali >>
rect 93 9732 157 9795
<< m1 >>
rect 93 9732 157 9795
<< viali >>
rect 100 9739 150 9788
<< locali >>
rect 1615 9732 1679 9795
<< m1 >>
rect 1615 9732 1679 9795
<< viali >>
rect 1622 9739 1672 9788
<< locali >>
rect 100 9118 1672 9167
<< locali >>
rect 93 9111 157 9174
<< m1 >>
rect 93 9111 157 9174
<< viali >>
rect 100 9118 150 9167
<< locali >>
rect 1615 9111 1679 9174
<< m1 >>
rect 1615 9111 1679 9174
<< viali >>
rect 1622 9118 1672 9167
<< locali >>
rect 100 11179 1672 11228
<< locali >>
rect 93 11172 157 11235
<< m1 >>
rect 93 11172 157 11235
<< viali >>
rect 100 11179 150 11228
<< locali >>
rect 1615 11172 1679 11235
<< m1 >>
rect 1615 11172 1679 11235
<< viali >>
rect 1622 11179 1672 11228
<< locali >>
rect 100 10558 1672 10607
<< locali >>
rect 93 10551 157 10614
<< m1 >>
rect 93 10551 157 10614
<< viali >>
rect 100 10558 150 10607
<< locali >>
rect 1615 10551 1679 10614
<< m1 >>
rect 1615 10551 1679 10614
<< viali >>
rect 1622 10558 1672 10607
<< locali >>
rect 100 10459 1672 10508
<< locali >>
rect 93 10452 157 10515
<< m1 >>
rect 93 10452 157 10515
<< viali >>
rect 100 10459 150 10508
<< locali >>
rect 1615 10452 1679 10515
<< m1 >>
rect 1615 10452 1679 10515
<< viali >>
rect 1622 10459 1672 10508
<< locali >>
rect 100 9838 1672 9887
<< locali >>
rect 93 9831 157 9894
<< m1 >>
rect 93 9831 157 9894
<< viali >>
rect 100 9838 150 9887
<< locali >>
rect 1615 9831 1679 9894
<< m1 >>
rect 1615 9831 1679 9894
<< viali >>
rect 1622 9838 1672 9887
<< locali >>
rect 100 13339 1672 13388
<< locali >>
rect 93 13332 157 13395
<< m1 >>
rect 93 13332 157 13395
<< viali >>
rect 100 13339 150 13388
<< locali >>
rect 1615 13332 1679 13395
<< m1 >>
rect 1615 13332 1679 13395
<< viali >>
rect 1622 13339 1672 13388
<< locali >>
rect 100 12718 1672 12767
<< locali >>
rect 93 12711 157 12774
<< m1 >>
rect 93 12711 157 12774
<< viali >>
rect 100 12718 150 12767
<< locali >>
rect 1615 12711 1679 12774
<< m1 >>
rect 1615 12711 1679 12774
<< viali >>
rect 1622 12718 1672 12767
<< locali >>
rect 100 8299 1672 8348
<< locali >>
rect 93 8292 157 8355
<< m1 >>
rect 93 8292 157 8355
<< viali >>
rect 100 8299 150 8348
<< locali >>
rect 1615 8292 1679 8355
<< m1 >>
rect 1615 8292 1679 8355
<< viali >>
rect 1622 8299 1672 8348
<< locali >>
rect 100 7678 1672 7727
<< locali >>
rect 93 7671 157 7734
<< m1 >>
rect 93 7671 157 7734
<< viali >>
rect 100 7678 150 7727
<< locali >>
rect 1615 7671 1679 7734
<< m1 >>
rect 1615 7671 1679 7734
<< viali >>
rect 1622 7678 1672 7727
<< locali >>
rect 100 12619 1672 12668
<< locali >>
rect 93 12612 157 12675
<< m1 >>
rect 93 12612 157 12675
<< viali >>
rect 100 12619 150 12668
<< locali >>
rect 1615 12612 1679 12675
<< m1 >>
rect 1615 12612 1679 12675
<< viali >>
rect 1622 12619 1672 12668
<< locali >>
rect 100 11998 1672 12047
<< locali >>
rect 93 11991 157 12054
<< m1 >>
rect 93 11991 157 12054
<< viali >>
rect 100 11998 150 12047
<< locali >>
rect 1615 11991 1679 12054
<< m1 >>
rect 1615 11991 1679 12054
<< viali >>
rect 1622 11998 1672 12047
<< locali >>
rect 100 9019 1672 9068
<< locali >>
rect 93 9012 157 9075
<< m1 >>
rect 93 9012 157 9075
<< viali >>
rect 100 9019 150 9068
<< locali >>
rect 1615 9012 1679 9075
<< m1 >>
rect 1615 9012 1679 9075
<< viali >>
rect 1622 9019 1672 9068
<< locali >>
rect 100 8398 1672 8447
<< locali >>
rect 93 8391 157 8454
<< m1 >>
rect 93 8391 157 8454
<< viali >>
rect 100 8398 150 8447
<< locali >>
rect 1615 8391 1679 8454
<< m1 >>
rect 1615 8391 1679 8454
<< viali >>
rect 1622 8398 1672 8447
<< locali >>
rect 100 11899 1672 11948
<< locali >>
rect 93 11892 157 11955
<< m1 >>
rect 93 11892 157 11955
<< viali >>
rect 100 11899 150 11948
<< locali >>
rect 1615 11892 1679 11955
<< m1 >>
rect 1615 11892 1679 11955
<< viali >>
rect 1622 11899 1672 11948
<< locali >>
rect 100 11278 1672 11327
<< locali >>
rect 93 11271 157 11334
<< m1 >>
rect 93 11271 157 11334
<< viali >>
rect 100 11278 150 11327
<< locali >>
rect 1615 11271 1679 11334
<< m1 >>
rect 1615 11271 1679 11334
<< viali >>
rect 1622 11278 1672 11327
<< locali >>
rect 0 3459 1772 3488
<< locali >>
rect 193 3452 787 3495
<< m1 >>
rect 193 3452 787 3495
<< m2 >>
rect 193 3452 787 3495
<< m3 >>
rect 193 3452 787 3495
<< viali >>
rect 200 3459 780 3488
<< via1 >>
rect 200 3459 780 3488
<< via2 >>
rect 200 3459 780 3488
<< locali >>
rect -7 3452 57 3495
<< m1 >>
rect -7 3452 57 3495
<< viali >>
rect 0 3459 50 3488
<< locali >>
rect 1715 3452 1779 3495
<< m1 >>
rect 1715 3452 1779 3495
<< viali >>
rect 1722 3459 1772 3488
use OTA U1_OTA 
transform 1 0 1822 0 1 0
box 0 0 2686 8956
<< labels >>
flabel locali s 0 14258 1772 14308 0 FreeSans 400 0 0 0 VDD
port 35 nsew signal bidirectional
flabel locali s 100 14158 1672 14208 0 FreeSans 400 0 0 0 VSS
port 36 nsew signal bidirectional
flabel m1 s 1204 1820 1300 1860 0 FreeSans 400 0 0 0 OUT
port 37 nsew signal bidirectional
<< properties >>
<< end >>