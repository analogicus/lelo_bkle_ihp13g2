magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747653241
<< checkpaint >>
rect 0 0 1 1
use LELOTR_NCHDL  None_MN2 ../LELO_TR_IHP13G2
timestamp 1747653241
transform 1 0 300 0 1 200
box 0 0 407 160
use LELOTR_NCHDL  None_MN3 ../LELO_TR_IHP13G2
timestamp 1747653241
transform 1 0 707 0 1 200
box 0 0 407 160
use LELOTR_PCHDL  None_MP2 ../LELO_TR_IHP13G2
timestamp 1747653241
transform 1 0 707 0 1 1080
box 0 0 407 160
use LELOTR_PCHDL  None_MP3 ../LELO_TR_IHP13G2
timestamp 1747653241
transform 1 0 300 0 1 1080
box 0 0 407 160
<< metal4 >>
rect 427 278 457 1029
<< metal3 >>
rect 427 999 985 1029
<< metal4 >>
rect 955 999 985 1158
<< metal3 >>
rect 420 992 464 1036
<< metal4 >>
rect 420 992 464 1036
<< via3 >>
rect 427 999 457 1029
<< metal3 >>
rect 948 992 992 1036
<< metal4 >>
rect 948 992 992 1036
<< via3 >>
rect 955 999 985 1029
<< metal4 >>
rect 830 278 860 917
<< metal3 >>
rect 542 887 860 917
<< metal4 >>
rect 542 887 572 1158
<< metal3 >>
rect 823 880 867 924
<< metal4 >>
rect 823 880 867 924
<< via3 >>
rect 830 887 860 917
<< metal3 >>
rect 535 880 579 924
<< metal4 >>
rect 535 880 579 924
<< via3 >>
rect 542 887 572 917
<< metal3 >>
rect 269 1101 412 1131
<< metal4 >>
rect 269 429 299 1131
<< metal3 >>
rect 269 429 1019 459
<< metal4 >>
rect 989 301 1019 459
<< metal4 >>
rect 989 301 1019 795
<< metal3 >>
rect 669 765 1019 795
<< metal4 >>
rect 669 765 699 1211
<< metal3 >>
rect 669 1181 812 1211
<< metal3 >>
rect 262 1094 306 1138
<< metal4 >>
rect 262 1094 306 1138
<< via3 >>
rect 269 1101 299 1131
<< metal3 >>
rect 262 422 306 466
<< metal4 >>
rect 262 422 306 466
<< via3 >>
rect 269 429 299 459
<< metal3 >>
rect 982 422 1026 466
<< metal4 >>
rect 982 422 1026 466
<< via3 >>
rect 989 429 1019 459
<< metal3 >>
rect 982 758 1026 802
<< metal4 >>
rect 982 758 1026 802
<< via3 >>
rect 989 765 1019 795
<< metal3 >>
rect 662 758 706 802
<< metal4 >>
rect 662 758 706 802
<< via3 >>
rect 669 765 699 795
<< metal3 >>
rect 662 1174 706 1218
<< metal4 >>
rect 662 1174 706 1218
<< via3 >>
rect 669 1181 699 1211
<< metal1 >>
rect 700 890 714 940
<< metal1 >>
rect 700 500 714 550
<< metal2 >>
rect 700 550 750 890
<< metal2 >>
rect 664 550 714 890
<< metal1 >>
rect 693 883 757 947
<< metal2 >>
rect 693 883 757 947
<< via1 >>
rect 700 890 750 940
<< metal1 >>
rect 693 493 757 557
<< metal2 >>
rect 693 493 757 557
<< via1 >>
rect 700 500 750 550
<< metal1 >>
rect 657 883 721 947
<< metal2 >>
rect 657 883 721 947
<< via1 >>
rect 664 890 714 940
<< metal1 >>
rect 657 493 721 557
<< metal2 >>
rect 657 493 721 557
<< via1 >>
rect 664 500 714 550
<< metal1 >>
rect 600 990 814 1040
<< metal1 >>
rect 600 400 814 450
<< metal2 >>
rect 600 450 650 990
<< metal2 >>
rect 764 450 814 990
<< metal1 >>
rect 593 983 657 1047
<< metal2 >>
rect 593 983 657 1047
<< via1 >>
rect 600 990 650 1040
<< metal1 >>
rect 593 393 657 457
<< metal2 >>
rect 593 393 657 457
<< via1 >>
rect 600 400 650 450
<< metal1 >>
rect 757 983 821 1047
<< metal2 >>
rect 757 983 821 1047
<< via1 >>
rect 764 990 814 1040
<< metal1 >>
rect 757 393 821 457
<< metal2 >>
rect 757 393 821 457
<< via1 >>
rect 764 400 814 450
<< metal1 >>
rect 392 263 494 297
<< metal2 >>
rect 392 263 494 297
<< metal3 >>
rect 392 263 494 297
<< metal4 >>
rect 392 263 494 297
<< via3 >>
rect 399 270 487 290
<< via2 >>
rect 399 270 487 290
<< via1 >>
rect 399 270 487 290
<< metal1 >>
rect 920 1143 1022 1177
<< metal2 >>
rect 920 1143 1022 1177
<< metal3 >>
rect 920 1143 1022 1177
<< metal4 >>
rect 920 1143 1022 1177
<< via3 >>
rect 927 1150 1015 1170
<< via2 >>
rect 927 1150 1015 1170
<< via1 >>
rect 927 1150 1015 1170
<< metal1 >>
rect 799 263 901 297
<< metal2 >>
rect 799 263 901 297
<< metal3 >>
rect 799 263 901 297
<< metal4 >>
rect 799 263 901 297
<< via3 >>
rect 806 270 894 290
<< via2 >>
rect 806 270 894 290
<< via1 >>
rect 806 270 894 290
<< metal1 >>
rect 513 1143 615 1177
<< metal2 >>
rect 513 1143 615 1177
<< metal3 >>
rect 513 1143 615 1177
<< metal4 >>
rect 513 1143 615 1177
<< via3 >>
rect 520 1150 608 1170
<< via2 >>
rect 520 1150 608 1170
<< via1 >>
rect 520 1150 608 1170
<< metal1 >>
rect 953 303 1055 337
<< metal2 >>
rect 953 303 1055 337
<< metal3 >>
rect 953 303 1055 337
<< metal4 >>
rect 953 303 1055 337
<< via3 >>
rect 960 310 1048 330
<< via2 >>
rect 960 310 1048 330
<< via1 >>
rect 960 310 1048 330
<< metal1 >>
rect 953 303 1055 337
<< metal2 >>
rect 953 303 1055 337
<< metal3 >>
rect 953 303 1055 337
<< metal4 >>
rect 953 303 1055 337
<< via3 >>
rect 960 310 1048 330
<< via2 >>
rect 960 310 1048 330
<< via1 >>
rect 960 310 1048 330
<< metal1 >>
rect 766 1183 868 1217
<< metal2 >>
rect 766 1183 868 1217
<< metal3 >>
rect 766 1183 868 1217
<< via2 >>
rect 773 1190 861 1210
<< via1 >>
rect 773 1190 861 1210
<< metal1 >>
rect 359 1103 461 1137
<< metal2 >>
rect 359 1103 461 1137
<< metal3 >>
rect 359 1103 461 1137
<< via2 >>
rect 366 1110 454 1130
<< via1 >>
rect 366 1110 454 1130
<< labels >>
flabel metal4 s 427 278 457 1029 0 FreeSans 400 0 0 0 A
port 23 nsew signal bidirectional
flabel metal4 s 830 278 860 917 0 FreeSans 400 0 0 0 B
port 24 nsew signal bidirectional
flabel metal3 s 269 1101 412 1131 0 FreeSans 400 0 0 0 Y
port 25 nsew signal bidirectional
flabel metal1 s 600 990 814 1040 0 FreeSans 400 0 0 0 AVDD
port 26 nsew signal bidirectional
flabel metal1 s 700 890 714 940 0 FreeSans 400 0 0 0 AVSS
port 27 nsew signal bidirectional
<< properties >>
<< end >>