magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747897834
<< checkpaint >>
rect 0 0 1 1
use LELOATR_NCH_4C5F0  diff1_MN1 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 1114
box 0 0 756 400
use LELOATR_NCH_4C5F0  diff1_MN2 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 1114
box 0 0 756 400
use LELOATR_PCH_4C5F0  load1_MP5 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 2614
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  load1_MP5_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 2374
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP6 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 2614
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  load1_MP6_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 2374
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP1 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 3014
box 0 0 756 400
use LELOATR_PCH_4C5F0  load1_MP2 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 3014
box 0 0 756 400
use LELOATR_NCH_4C5F0  mirror2_MN4 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 1514
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN4_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 1914
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN3 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 1514
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN3_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 1914
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror1_MN5 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 714
box 0 0 756 400
use LELOATR_NCH_4CTAPBOT  mirror1_MN5_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 474
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror1_MN6 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 714
box 0 0 756 400
use LELOATR_NCH_4CTAPBOT  mirror1_MN6_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 474
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP3 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 3414
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP3_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 738 0 1 3814
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP4 ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 3414
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP4_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1747897834
transform 1 0 1494 0 1 3814
box 0 0 756 240
<< metal3 >>
rect 1998 2635 2157 2665
<< metal4 >>
rect 2127 731 2157 2665
<< metal3 >>
rect 1998 731 2157 761
<< metal3 >>
rect 2120 2628 2164 2672
<< metal4 >>
rect 2120 2628 2164 2672
<< via3 >>
rect 2127 2635 2157 2665
<< metal3 >>
rect 2120 724 2164 768
<< metal4 >>
rect 2120 724 2164 768
<< via3 >>
rect 2127 731 2157 761
<< metal3 >>
rect 863 1693 1615 1723
<< metal4 >>
rect 1605 3213 1635 3628
<< metal4 >>
rect 1605 3438 1635 3628
<< metal3 >>
rect 1221 3438 1635 3468
<< metal3 >>
rect 853 3438 1251 3468
<< metal4 >>
rect 853 3198 883 3468
<< metal3 >>
rect 725 3198 883 3228
<< metal4 >>
rect 725 1134 755 3228
<< metal3 >>
rect 725 1134 1236 1164
<< metal3 >>
rect 1598 3431 1642 3475
<< metal4 >>
rect 1598 3431 1642 3475
<< via3 >>
rect 1605 3438 1635 3468
<< metal3 >>
rect 846 3431 890 3475
<< metal4 >>
rect 846 3431 890 3475
<< via3 >>
rect 853 3438 883 3468
<< metal3 >>
rect 846 3191 890 3235
<< metal4 >>
rect 846 3191 890 3235
<< via3 >>
rect 853 3198 883 3228
<< metal3 >>
rect 718 3191 762 3235
<< metal4 >>
rect 718 3191 762 3235
<< via3 >>
rect 725 3198 755 3228
<< metal3 >>
rect 718 1127 762 1171
<< metal4 >>
rect 718 1127 762 1171
<< via3 >>
rect 725 1134 755 1164
<< metal4 >>
rect 1216 1290 1246 1545
<< metal3 >>
rect 976 1290 1246 1320
<< metal4 >>
rect 976 1290 1006 1448
<< metal3 >>
rect 976 1418 1262 1448
<< metal3 >>
rect 1232 1418 1743 1448
<< metal3 >>
rect 1209 1283 1253 1327
<< metal4 >>
rect 1209 1283 1253 1327
<< via3 >>
rect 1216 1290 1246 1320
<< metal3 >>
rect 969 1283 1013 1327
<< metal4 >>
rect 969 1283 1013 1327
<< via3 >>
rect 976 1290 1006 1320
<< metal3 >>
rect 969 1411 1013 1455
<< metal4 >>
rect 969 1411 1013 1455
<< via3 >>
rect 976 1418 1006 1448
<< metal3 >>
rect 625 3598 864 3628
<< metal4 >>
rect 625 2798 655 3628
<< metal3 >>
rect 625 2798 879 2828
<< metal3 >>
rect 849 2798 1631 2828
<< metal4 >>
rect 1601 2798 1631 3052
<< metal3 >>
rect 1601 3022 1871 3052
<< metal4 >>
rect 1841 3022 1871 3180
<< metal3 >>
rect 1841 3150 2015 3180
<< metal4 >>
rect 1985 3150 2015 3468
<< metal3 >>
rect 1985 3438 2255 3468
<< metal4 >>
rect 2225 1134 2255 3468
<< metal3 >>
rect 2000 1134 2255 1164
<< metal3 >>
rect 618 3591 662 3635
<< metal4 >>
rect 618 3591 662 3635
<< via3 >>
rect 625 3598 655 3628
<< metal3 >>
rect 618 2791 662 2835
<< metal4 >>
rect 618 2791 662 2835
<< via3 >>
rect 625 2798 655 2828
<< metal3 >>
rect 1594 2791 1638 2835
<< metal4 >>
rect 1594 2791 1638 2835
<< via3 >>
rect 1601 2798 1631 2828
<< metal3 >>
rect 1594 3015 1638 3059
<< metal4 >>
rect 1594 3015 1638 3059
<< via3 >>
rect 1601 3022 1631 3052
<< metal3 >>
rect 1834 3015 1878 3059
<< metal4 >>
rect 1834 3015 1878 3059
<< via3 >>
rect 1841 3022 1871 3052
<< metal3 >>
rect 1834 3143 1878 3187
<< metal4 >>
rect 1834 3143 1878 3187
<< via3 >>
rect 1841 3150 1871 3180
<< metal3 >>
rect 1978 3143 2022 3187
<< metal4 >>
rect 1978 3143 2022 3187
<< via3 >>
rect 1985 3150 2015 3180
<< metal3 >>
rect 1978 3431 2022 3475
<< metal4 >>
rect 1978 3431 2022 3475
<< via3 >>
rect 1985 3438 2015 3468
<< metal3 >>
rect 2218 3431 2262 3475
<< metal4 >>
rect 2218 3431 2262 3475
<< via3 >>
rect 2225 3438 2255 3468
<< metal3 >>
rect 2218 1127 2262 1171
<< metal4 >>
rect 2218 1127 2262 1171
<< via3 >>
rect 2225 1134 2255 1164
<< metal3 >>
rect 852 894 1619 924
<< metal3 >>
rect 852 894 1394 924
<< metal4 >>
rect 1364 894 1394 3068
<< metal3 >>
rect 1235 3038 1394 3068
<< metal3 >>
rect 1357 887 1401 931
<< metal4 >>
rect 1357 887 1401 931
<< via3 >>
rect 1364 894 1394 924
<< metal3 >>
rect 1357 3031 1401 3075
<< metal4 >>
rect 1357 3031 1401 3075
<< via3 >>
rect 1364 3038 1394 3068
<< metal1 >>
rect 100 4378 2888 4428
<< metal1 >>
rect 100 100 2888 150
<< metal2 >>
rect 100 150 150 4378
<< metal2 >>
rect 2838 150 2888 4378
<< metal1 >>
rect 93 4371 157 4435
<< metal2 >>
rect 93 4371 157 4435
<< via1 >>
rect 100 4378 150 4428
<< metal1 >>
rect 93 93 157 157
<< metal2 >>
rect 93 93 157 157
<< via1 >>
rect 100 100 150 150
<< metal1 >>
rect 2831 4371 2895 4435
<< metal2 >>
rect 2831 4371 2895 4435
<< via1 >>
rect 2838 4378 2888 4428
<< metal1 >>
rect 2831 93 2895 157
<< metal2 >>
rect 2831 93 2895 157
<< via1 >>
rect 2838 100 2888 150
<< metal1 >>
rect 0 4478 2988 4528
<< metal1 >>
rect 0 0 2988 50
<< metal2 >>
rect 0 50 50 4478
<< metal2 >>
rect 2938 50 2988 4478
<< metal1 >>
rect -7 4471 57 4535
<< metal2 >>
rect -7 4471 57 4535
<< via1 >>
rect 0 4478 50 4528
<< metal1 >>
rect -7 -7 57 57
<< metal2 >>
rect -7 -7 57 57
<< via1 >>
rect 0 0 50 50
<< metal1 >>
rect 2931 4471 2995 4535
<< metal2 >>
rect 2931 4471 2995 4535
<< via1 >>
rect 2938 4478 2988 4528
<< metal1 >>
rect 2931 -7 2995 57
<< metal2 >>
rect 2931 -7 2995 57
<< via1 >>
rect 2938 0 2988 50
<< metal1 >>
rect 675 2914 1053 2954
<< metal1 >>
rect 1179 2794 1389 2834
<< metal1 >>
rect 1431 2914 1809 2954
<< metal1 >>
rect 675 3314 1053 3354
<< metal1 >>
rect 1431 3314 1809 3354
<< metal1 >>
rect 1935 3194 2145 3234
<< metal1 >>
rect 675 1814 1053 1854
<< metal1 >>
rect 1431 1814 1809 1854
<< metal1 >>
rect 1935 1694 2145 1734
<< metal1 >>
rect 675 1014 1053 1054
<< metal1 >>
rect 1179 894 1389 934
<< metal1 >>
rect 1431 1014 1809 1054
<< metal1 >>
rect 675 3714 1053 3754
<< metal1 >>
rect 1431 3714 1809 3754
<< metal1 >>
rect 0 2431 2988 2557
<< metal1 >>
rect -7 2424 57 2564
<< metal2 >>
rect -7 2424 57 2564
<< via1 >>
rect 0 2431 50 2557
<< metal1 >>
rect 2931 2424 2995 2564
<< metal2 >>
rect 2931 2424 2995 2564
<< via1 >>
rect 2938 2431 2988 2557
<< metal1 >>
rect 100 1971 2888 2097
<< metal1 >>
rect 93 1964 157 2104
<< metal2 >>
rect 93 1964 157 2104
<< via1 >>
rect 100 1971 150 2097
<< metal1 >>
rect 2831 1964 2895 2104
<< metal2 >>
rect 2831 1964 2895 2104
<< via1 >>
rect 2838 1971 2888 2097
<< metal1 >>
rect 100 531 2888 657
<< metal1 >>
rect 93 524 157 664
<< metal2 >>
rect 93 524 157 664
<< via1 >>
rect 100 531 150 657
<< metal1 >>
rect 2831 524 2895 664
<< metal2 >>
rect 2831 524 2895 664
<< via1 >>
rect 2838 531 2888 657
<< metal1 >>
rect 0 3871 2988 3997
<< metal1 >>
rect -7 3864 57 4004
<< metal2 >>
rect -7 3864 57 4004
<< via1 >>
rect 0 3871 50 3997
<< metal1 >>
rect 2931 3864 2995 4004
<< metal2 >>
rect 2931 3864 2995 4004
<< via1 >>
rect 2938 3871 2988 3997
<< metal2 >>
rect 1928 2627 2068 2681
<< metal3 >>
rect 1928 2627 2068 2681
<< via2 >>
rect 1935 2634 2061 2674
<< metal2 >>
rect 1928 727 2068 781
<< metal3 >>
rect 1928 727 2068 781
<< via2 >>
rect 1935 734 2061 774
<< metal2 >>
rect 836 1687 892 1741
<< metal3 >>
rect 836 1687 892 1741
<< via2 >>
rect 843 1694 885 1734
<< metal2 >>
rect 1592 1687 1648 1741
<< metal3 >>
rect 1592 1687 1648 1741
<< via2 >>
rect 1599 1694 1641 1734
<< metal2 >>
rect 1172 1127 1312 1181
<< metal3 >>
rect 1172 1127 1312 1181
<< via2 >>
rect 1179 1134 1305 1174
<< metal2 >>
rect 836 3187 892 3241
<< metal3 >>
rect 836 3187 892 3241
<< metal4 >>
rect 836 3187 892 3241
<< via3 >>
rect 843 3194 885 3234
<< via2 >>
rect 843 3194 885 3234
<< metal2 >>
rect 836 3187 892 3241
<< metal3 >>
rect 836 3187 892 3241
<< via2 >>
rect 843 3194 885 3234
<< metal2 >>
rect 1592 3187 1648 3241
<< metal3 >>
rect 1592 3187 1648 3241
<< metal4 >>
rect 1592 3187 1648 3241
<< via3 >>
rect 1599 3194 1641 3234
<< via2 >>
rect 1599 3194 1641 3234
<< metal2 >>
rect 1172 3427 1312 3481
<< metal3 >>
rect 1172 3427 1312 3481
<< via2 >>
rect 1179 3434 1305 3474
<< metal2 >>
rect 1172 3427 1312 3481
<< metal3 >>
rect 1172 3427 1312 3481
<< via2 >>
rect 1179 3434 1305 3474
<< metal2 >>
rect 1592 3587 1648 3641
<< metal3 >>
rect 1592 3587 1648 3641
<< metal4 >>
rect 1592 3587 1648 3641
<< via3 >>
rect 1599 3594 1641 3634
<< via2 >>
rect 1599 3594 1641 3634
<< metal2 >>
rect 1592 3587 1648 3641
<< metal3 >>
rect 1592 3587 1648 3641
<< metal4 >>
rect 1592 3587 1648 3641
<< via3 >>
rect 1599 3594 1641 3634
<< via2 >>
rect 1599 3594 1641 3634
<< metal2 >>
rect 920 1407 1060 1461
<< metal3 >>
rect 920 1407 1060 1461
<< metal4 >>
rect 920 1407 1060 1461
<< via3 >>
rect 927 1414 1053 1454
<< via2 >>
rect 927 1414 1053 1454
<< metal2 >>
rect 920 1407 1060 1461
<< metal3 >>
rect 920 1407 1060 1461
<< via2 >>
rect 927 1414 1053 1454
<< metal2 >>
rect 1676 1407 1816 1461
<< metal3 >>
rect 1676 1407 1816 1461
<< via2 >>
rect 1683 1414 1809 1454
<< metal2 >>
rect 1172 1527 1312 1581
<< metal3 >>
rect 1172 1527 1312 1581
<< metal4 >>
rect 1172 1527 1312 1581
<< via3 >>
rect 1179 1534 1305 1574
<< via2 >>
rect 1179 1534 1305 1574
<< metal2 >>
rect 1928 1127 2068 1181
<< metal3 >>
rect 1928 1127 2068 1181
<< via2 >>
rect 1935 1134 2061 1174
<< metal2 >>
rect 836 2787 892 2841
<< metal3 >>
rect 836 2787 892 2841
<< via2 >>
rect 843 2794 885 2834
<< metal2 >>
rect 836 2787 892 2841
<< metal3 >>
rect 836 2787 892 2841
<< via2 >>
rect 843 2794 885 2834
<< metal2 >>
rect 1592 2787 1648 2841
<< metal3 >>
rect 1592 2787 1648 2841
<< via2 >>
rect 1599 2794 1641 2834
<< metal2 >>
rect 1592 2787 1648 2841
<< metal3 >>
rect 1592 2787 1648 2841
<< metal4 >>
rect 1592 2787 1648 2841
<< via3 >>
rect 1599 2794 1641 2834
<< via2 >>
rect 1599 2794 1641 2834
<< metal2 >>
rect 836 3587 892 3641
<< metal3 >>
rect 836 3587 892 3641
<< via2 >>
rect 843 3594 885 3634
<< metal2 >>
rect 1928 3427 2068 3481
<< metal3 >>
rect 1928 3427 2068 3481
<< metal4 >>
rect 1928 3427 2068 3481
<< via3 >>
rect 1935 3434 2061 3474
<< via2 >>
rect 1935 3434 2061 3474
<< metal2 >>
rect 1928 3427 2068 3481
<< metal3 >>
rect 1928 3427 2068 3481
<< via2 >>
rect 1935 3434 2061 3474
<< metal2 >>
rect 1172 3027 1312 3081
<< metal3 >>
rect 1172 3027 1312 3081
<< via2 >>
rect 1179 3034 1305 3074
<< metal2 >>
rect 836 887 892 941
<< metal3 >>
rect 836 887 892 941
<< via2 >>
rect 843 894 885 934
<< metal2 >>
rect 836 887 892 941
<< metal3 >>
rect 836 887 892 941
<< via2 >>
rect 843 894 885 934
<< metal2 >>
rect 1592 887 1648 941
<< metal3 >>
rect 1592 887 1648 941
<< via2 >>
rect 1599 894 1641 934
<< labels >>
flabel metal1 s 100 4378 2888 4428 0 FreeSans 400 0 0 0 VSS
port 4 nsew signal bidirectional
flabel metal1 s 0 4478 2988 4528 0 FreeSans 400 0 0 0 VDD
port 5 nsew signal bidirectional
flabel metal2 s 843 1294 885 1334 0 FreeSans 400 0 0 0 VIP
port 6 nsew signal bidirectional
flabel metal2 s 1599 1294 1641 1334 0 FreeSans 400 0 0 0 VIN
port 7 nsew signal bidirectional
flabel metal3 s 1998 2635 2157 2665 0 FreeSans 400 0 0 0 VO
port 8 nsew signal bidirectional
flabel metal3 s 863 1693 1615 1723 0 FreeSans 400 0 0 0 I_BIAS
port 9 nsew signal bidirectional
<< properties >>
<< end >>