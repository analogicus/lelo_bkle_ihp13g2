magic
tech ihp-sg13g2
magscale 1 1
timestamp 1748119001
<< checkpaint >>
rect 0 0 1 1
use LELOATR_NCH_4C5F0  diff1_MN1 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 2002
box 0 0 756 400
use LELOATR_NCH_4CTAPBOT  diff1_MN1_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 1762
box 0 0 756 240
use LELOATR_NCH_4C5F0  diff1_MN2 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 2002
box 0 0 756 400
use LELOATR_NCH_4CTAPBOT  diff1_MN2_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 1762
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP5 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 902
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP5_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 1302
box 0 0 756 240
use LELOATR_PCH_4CTAPBOT  load1_MP5_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 662
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP6 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 902
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP6_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 1302
box 0 0 756 240
use LELOATR_PCH_4CTAPBOT  load1_MP6_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 662
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP1 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 502
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  load1_MP1_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 262
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP2 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 502
box 0 0 756 400
use LELOATR_PCH_4CTAPBOT  load1_MP2_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 262
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN4 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 2402
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN4_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 2802
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror2_MN3 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 2402
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror2_MN3_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 2802
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror1_MN5 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 2402
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror1_MN5_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 2802
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror1_MN5_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 2573 0 1 2162
box 0 0 756 240
use LELOATR_NCH_4C5F0  mirror1_MN6 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 2402
box 0 0 756 400
use LELOATR_NCH_4CTAPTOP  mirror1_MN6_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 2802
box 0 0 756 240
use LELOATR_NCH_4CTAPBOT  mirror1_MN6_TAPBOT ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 305 0 1 2162
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP3 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 902
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP3_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1817 0 1 1302
box 0 0 756 240
use LELOATR_PCH_4C5F0  load1_MP4 ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 902
box 0 0 756 400
use LELOATR_PCH_4CTAPTOP  load1_MP4_TAPTOP ../LELO_ATR_IHP13G2
timestamp 1748119001
transform 1 0 1061 0 1 1302
box 0 0 756 240
<< metal4 >>
rect 788 936 818 2440
<< metal3 >>
rect 1184 2583 1936 2613
<< metal4 >>
rect 1171 684 1201 1099
<< metal3 >>
rect 1171 684 1953 714
<< metal3 >>
rect 1923 684 2337 714
<< metal4 >>
rect 2307 684 2337 954
<< metal4 >>
rect 2307 924 2337 2043
<< metal3 >>
rect 1164 677 1208 721
<< metal4 >>
rect 1164 677 1208 721
<< via3 >>
rect 1171 684 1201 714
<< metal3 >>
rect 2300 677 2344 721
<< metal4 >>
rect 2300 677 2344 721
<< via3 >>
rect 2307 684 2337 714
<< metal4 >>
rect 1554 2179 1584 2434
<< metal3 >>
rect 1298 2179 1584 2209
<< metal4 >>
rect 1298 2179 1328 2337
<< metal3 >>
rect 1298 2307 1600 2337
<< metal3 >>
rect 1570 2307 2065 2337
<< metal3 >>
rect 1547 2172 1591 2216
<< metal4 >>
rect 1547 2172 1591 2216
<< via3 >>
rect 1554 2179 1584 2209
<< metal3 >>
rect 1291 2172 1335 2216
<< metal4 >>
rect 1291 2172 1335 2216
<< via3 >>
rect 1298 2179 1328 2209
<< metal3 >>
rect 1291 2300 1335 2344
<< metal4 >>
rect 1291 2300 1335 2344
<< via3 >>
rect 1298 2307 1328 2337
<< metal3 >>
rect 434 1084 1025 1114
<< metal4 >>
rect 995 924 1025 1114
<< metal3 >>
rect 995 924 1585 954
<< metal4 >>
rect 1555 924 1585 2058
<< metal4 >>
rect 1555 1084 1585 2058
<< metal3 >>
rect 1555 1084 1953 1114
<< metal3 >>
rect 1923 1084 2690 1114
<< metal3 >>
rect 988 1077 1032 1121
<< metal4 >>
rect 988 1077 1032 1121
<< via3 >>
rect 995 1084 1025 1114
<< metal3 >>
rect 988 917 1032 961
<< metal4 >>
rect 988 917 1032 961
<< via3 >>
rect 995 924 1025 954
<< metal3 >>
rect 1548 917 1592 961
<< metal4 >>
rect 1548 917 1592 961
<< via3 >>
rect 1555 924 1585 954
<< metal3 >>
rect 1548 1077 1592 1121
<< metal4 >>
rect 1548 1077 1592 1121
<< via3 >>
rect 1555 1084 1585 1114
<< metal4 >>
rect 419 2601 449 2824
<< metal3 >>
rect 419 2794 2705 2824
<< metal4 >>
rect 2675 2586 2705 2824
<< metal4 >>
rect 2675 1322 2705 2616
<< metal3 >>
rect 1715 1322 2705 1352
<< metal4 >>
rect 1715 522 1745 1352
<< metal3 >>
rect 1570 522 1745 552
<< metal3 >>
rect 412 2787 456 2831
<< metal4 >>
rect 412 2787 456 2831
<< via3 >>
rect 419 2794 449 2824
<< metal3 >>
rect 2668 2787 2712 2831
<< metal4 >>
rect 2668 2787 2712 2831
<< via3 >>
rect 2675 2794 2705 2824
<< metal3 >>
rect 2668 1315 2712 1359
<< metal4 >>
rect 2668 1315 2712 1359
<< via3 >>
rect 2675 1322 2705 1352
<< metal3 >>
rect 1708 1315 1752 1359
<< metal4 >>
rect 1708 1315 1752 1359
<< via3 >>
rect 1715 1322 1745 1352
<< metal3 >>
rect 1708 515 1752 559
<< metal4 >>
rect 1708 515 1752 559
<< via3 >>
rect 1715 522 1745 552
<< metal1 >>
rect 100 3154 3534 3204
<< metal1 >>
rect 100 100 3534 150
<< metal2 >>
rect 100 150 150 3154
<< metal2 >>
rect 3484 150 3534 3154
<< metal1 >>
rect 93 3147 157 3211
<< metal2 >>
rect 93 3147 157 3211
<< via1 >>
rect 100 3154 150 3204
<< metal1 >>
rect 93 93 157 157
<< metal2 >>
rect 93 93 157 157
<< via1 >>
rect 100 100 150 150
<< metal1 >>
rect 3477 3147 3541 3211
<< metal2 >>
rect 3477 3147 3541 3211
<< via1 >>
rect 3484 3154 3534 3204
<< metal1 >>
rect 3477 93 3541 157
<< metal2 >>
rect 3477 93 3541 157
<< via1 >>
rect 3484 100 3534 150
<< metal1 >>
rect 0 3254 3634 3304
<< metal1 >>
rect 0 0 3634 50
<< metal2 >>
rect 0 50 50 3254
<< metal2 >>
rect 3584 50 3634 3254
<< metal1 >>
rect -7 3247 57 3311
<< metal2 >>
rect -7 3247 57 3311
<< via1 >>
rect 0 3254 50 3304
<< metal1 >>
rect -7 -7 57 57
<< metal2 >>
rect -7 -7 57 57
<< via1 >>
rect 0 0 50 50
<< metal1 >>
rect 3577 3247 3641 3311
<< metal2 >>
rect 3577 3247 3641 3311
<< via1 >>
rect 3584 3254 3634 3304
<< metal1 >>
rect 3577 -7 3641 57
<< metal2 >>
rect 3577 -7 3641 57
<< via1 >>
rect 3584 0 3634 50
<< metal1 >>
rect 2510 1202 2888 1242
<< metal1 >>
rect 3014 1082 3224 1122
<< metal1 >>
rect 242 1202 620 1242
<< metal1 >>
rect 998 802 1376 842
<< metal1 >>
rect 1754 802 2132 842
<< metal1 >>
rect 2258 682 2468 722
<< metal1 >>
rect 998 2702 1376 2742
<< metal1 >>
rect 1754 2702 2132 2742
<< metal1 >>
rect 2258 2582 2468 2622
<< metal1 >>
rect 2510 2702 2888 2742
<< metal1 >>
rect 3014 2582 3224 2622
<< metal1 >>
rect 242 2702 620 2742
<< metal1 >>
rect 1754 1202 2132 1242
<< metal1 >>
rect 998 1202 1376 1242
<< metal1 >>
rect 100 1819 3534 1945
<< metal1 >>
rect 93 1812 157 1952
<< metal2 >>
rect 93 1812 157 1952
<< via1 >>
rect 100 1819 150 1945
<< metal1 >>
rect 3477 1812 3541 1952
<< metal2 >>
rect 3477 1812 3541 1952
<< via1 >>
rect 3484 1819 3534 1945
<< metal1 >>
rect 0 1359 3634 1485
<< metal1 >>
rect -7 1352 57 1492
<< metal2 >>
rect -7 1352 57 1492
<< via1 >>
rect 0 1359 50 1485
<< metal1 >>
rect 3577 1352 3641 1492
<< metal2 >>
rect 3577 1352 3641 1492
<< via1 >>
rect 3584 1359 3634 1485
<< metal1 >>
rect 0 319 3634 445
<< metal1 >>
rect -7 312 57 452
<< metal2 >>
rect -7 312 57 452
<< via1 >>
rect 0 319 50 445
<< metal1 >>
rect 3577 312 3641 452
<< metal2 >>
rect 3577 312 3641 452
<< via1 >>
rect 3584 319 3634 445
<< metal1 >>
rect 100 2859 3534 2985
<< metal1 >>
rect 93 2852 157 2992
<< metal2 >>
rect 93 2852 157 2992
<< via1 >>
rect 100 2859 150 2985
<< metal1 >>
rect 3477 2852 3541 2992
<< metal2 >>
rect 3477 2852 3541 2992
<< via1 >>
rect 3484 2859 3534 2985
<< metal2 >>
rect 739 915 879 969
<< metal3 >>
rect 739 915 879 969
<< metal4 >>
rect 739 915 879 969
<< via3 >>
rect 746 922 872 962
<< via2 >>
rect 746 922 872 962
<< metal2 >>
rect 739 2415 879 2469
<< metal3 >>
rect 739 2415 879 2469
<< metal4 >>
rect 739 2415 879 2469
<< via3 >>
rect 746 2422 872 2462
<< via2 >>
rect 746 2422 872 2462
<< metal2 >>
rect 1159 2575 1215 2629
<< metal3 >>
rect 1159 2575 1215 2629
<< via2 >>
rect 1166 2582 1208 2622
<< metal2 >>
rect 1915 2575 1971 2629
<< metal3 >>
rect 1915 2575 1971 2629
<< via2 >>
rect 1922 2582 1964 2622
<< metal2 >>
rect 2251 2015 2391 2069
<< metal3 >>
rect 2251 2015 2391 2069
<< metal4 >>
rect 2251 2015 2391 2069
<< via3 >>
rect 2258 2022 2384 2062
<< via2 >>
rect 2258 2022 2384 2062
<< metal2 >>
rect 1159 675 1215 729
<< metal3 >>
rect 1159 675 1215 729
<< metal4 >>
rect 1159 675 1215 729
<< via3 >>
rect 1166 682 1208 722
<< via2 >>
rect 1166 682 1208 722
<< metal2 >>
rect 1159 675 1215 729
<< metal3 >>
rect 1159 675 1215 729
<< via2 >>
rect 1166 682 1208 722
<< metal2 >>
rect 1915 675 1971 729
<< metal3 >>
rect 1915 675 1971 729
<< via2 >>
rect 1922 682 1964 722
<< metal2 >>
rect 1915 675 1971 729
<< metal3 >>
rect 1915 675 1971 729
<< via2 >>
rect 1922 682 1964 722
<< metal2 >>
rect 2251 915 2391 969
<< metal3 >>
rect 2251 915 2391 969
<< metal4 >>
rect 2251 915 2391 969
<< via3 >>
rect 2258 922 2384 962
<< via2 >>
rect 2258 922 2384 962
<< metal2 >>
rect 2251 915 2391 969
<< metal3 >>
rect 2251 915 2391 969
<< metal4 >>
rect 2251 915 2391 969
<< via3 >>
rect 2258 922 2384 962
<< via2 >>
rect 2258 922 2384 962
<< metal2 >>
rect 1159 1075 1215 1129
<< metal3 >>
rect 1159 1075 1215 1129
<< metal4 >>
rect 1159 1075 1215 1129
<< via3 >>
rect 1166 1082 1208 1122
<< via2 >>
rect 1166 1082 1208 1122
<< metal2 >>
rect 1999 2295 2139 2349
<< metal3 >>
rect 1999 2295 2139 2349
<< via2 >>
rect 2006 2302 2132 2342
<< metal2 >>
rect 1243 2295 1383 2349
<< metal3 >>
rect 1243 2295 1383 2349
<< metal4 >>
rect 1243 2295 1383 2349
<< via3 >>
rect 1250 2302 1376 2342
<< via2 >>
rect 1250 2302 1376 2342
<< metal2 >>
rect 1243 2295 1383 2349
<< metal3 >>
rect 1243 2295 1383 2349
<< via2 >>
rect 1250 2302 1376 2342
<< metal2 >>
rect 1495 2415 1635 2469
<< metal3 >>
rect 1495 2415 1635 2469
<< metal4 >>
rect 1495 2415 1635 2469
<< via3 >>
rect 1502 2422 1628 2462
<< via2 >>
rect 1502 2422 1628 2462
<< metal2 >>
rect 1495 2015 1635 2069
<< metal3 >>
rect 1495 2015 1635 2069
<< metal4 >>
rect 1495 2015 1635 2069
<< via3 >>
rect 1502 2022 1628 2062
<< via2 >>
rect 1502 2022 1628 2062
<< metal2 >>
rect 1495 2015 1635 2069
<< metal3 >>
rect 1495 2015 1635 2069
<< metal4 >>
rect 1495 2015 1635 2069
<< via3 >>
rect 1502 2022 1628 2062
<< via2 >>
rect 1502 2022 1628 2062
<< metal2 >>
rect 2671 1075 2727 1129
<< metal3 >>
rect 2671 1075 2727 1129
<< via2 >>
rect 2678 1082 2720 1122
<< metal2 >>
rect 403 1075 459 1129
<< metal3 >>
rect 403 1075 459 1129
<< via2 >>
rect 410 1082 452 1122
<< metal2 >>
rect 1915 1075 1971 1129
<< metal3 >>
rect 1915 1075 1971 1129
<< via2 >>
rect 1922 1082 1964 1122
<< metal2 >>
rect 1915 1075 1971 1129
<< metal3 >>
rect 1915 1075 1971 1129
<< via2 >>
rect 1922 1082 1964 1122
<< metal2 >>
rect 1495 915 1635 969
<< metal3 >>
rect 1495 915 1635 969
<< via2 >>
rect 1502 922 1628 962
<< metal2 >>
rect 1495 915 1635 969
<< metal3 >>
rect 1495 915 1635 969
<< metal4 >>
rect 1495 915 1635 969
<< via3 >>
rect 1502 922 1628 962
<< via2 >>
rect 1502 922 1628 962
<< metal2 >>
rect 1495 515 1635 569
<< metal3 >>
rect 1495 515 1635 569
<< via2 >>
rect 1502 522 1628 562
<< metal2 >>
rect 2671 2575 2727 2629
<< metal3 >>
rect 2671 2575 2727 2629
<< metal4 >>
rect 2671 2575 2727 2629
<< via3 >>
rect 2678 2582 2720 2622
<< via2 >>
rect 2678 2582 2720 2622
<< metal2 >>
rect 2671 2575 2727 2629
<< metal3 >>
rect 2671 2575 2727 2629
<< metal4 >>
rect 2671 2575 2727 2629
<< via3 >>
rect 2678 2582 2720 2622
<< via2 >>
rect 2678 2582 2720 2622
<< metal2 >>
rect 403 2575 459 2629
<< metal3 >>
rect 403 2575 459 2629
<< metal4 >>
rect 403 2575 459 2629
<< via3 >>
rect 410 2582 452 2622
<< via2 >>
rect 410 2582 452 2622
<< labels >>
flabel metal1 s 100 3154 3534 3204 0 FreeSans 400 0 0 0 VSS
port 4 nsew signal bidirectional
flabel metal1 s 0 3254 3634 3304 0 FreeSans 400 0 0 0 VDD
port 5 nsew signal bidirectional
flabel metal2 s 1922 2182 1964 2222 0 FreeSans 400 0 0 0 VIP
port 6 nsew signal bidirectional
flabel metal2 s 1166 2182 1208 2222 0 FreeSans 400 0 0 0 VIN
port 7 nsew signal bidirectional
flabel metal4 s 788 936 818 2440 0 FreeSans 400 0 0 0 VO
port 8 nsew signal bidirectional
flabel metal3 s 1184 2583 1936 2613 0 FreeSans 400 0 0 0 I_BIAS
port 9 nsew signal bidirectional
<< properties >>
<< end >>