magic
tech ihp-sg13g2
magscale 1 1
timestamp 1747994531
<< checkpaint >>
rect 0 0 1 1
<< metal1 >>
rect -100 4030 5765 4080
<< metal1 >>
rect -100 -100 5765 -50
<< metal2 >>
rect -100 -50 -50 4030
<< metal2 >>
rect 5715 -50 5765 4030
<< metal1 >>
rect -107 4023 -43 4087
<< metal2 >>
rect -107 4023 -43 4087
<< via1 >>
rect -100 4030 -50 4080
<< metal1 >>
rect -107 -107 -43 -43
<< metal2 >>
rect -107 -107 -43 -43
<< via1 >>
rect -100 -100 -50 -50
<< metal1 >>
rect 5708 4023 5772 4087
<< metal2 >>
rect 5708 4023 5772 4087
<< via1 >>
rect 5715 4030 5765 4080
<< metal1 >>
rect 5708 -107 5772 -43
<< metal2 >>
rect 5708 -107 5772 -43
<< via1 >>
rect 5715 -100 5765 -50
<< metal1 >>
rect -200 4130 5865 4180
<< metal1 >>
rect -200 -200 5865 -150
<< metal2 >>
rect -200 -150 -150 4130
<< metal2 >>
rect 5815 -150 5865 4130
<< metal1 >>
rect -207 4123 -143 4187
<< metal2 >>
rect -207 4123 -143 4187
<< via1 >>
rect -200 4130 -150 4180
<< metal1 >>
rect -207 -207 -143 -143
<< metal2 >>
rect -207 -207 -143 -143
<< via1 >>
rect -200 -200 -150 -150
<< metal1 >>
rect 5808 4123 5872 4187
<< metal2 >>
rect 5808 4123 5872 4187
<< via1 >>
rect 5815 4130 5865 4180
<< metal1 >>
rect 5808 -207 5872 -143
<< metal2 >>
rect 5808 -207 5872 -143
<< via1 >>
rect 5815 -200 5865 -150
use OTA U1_OTA 
transform 1 0 0 0 1 0
box 0 0 5715 4030
<< labels >>
flabel metal1 s -200 4130 5865 4180 0 FreeSans 400 0 0 0 VDD_1V8
port 51 nsew signal bidirectional
flabel metal1 s -100 4030 5765 4080 0 FreeSans 400 0 0 0 VSS
port 52 nsew signal bidirectional
<< properties >>
<< end >>